library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity turkey_shoot_bank_c is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of turkey_shoot_bank_c is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"28",X"43",X"29",X"20",X"31",X"39",
		X"38",X"34",X"2C",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",
		X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"00",X"0C",X"CC",
		X"C0",X"00",X"00",X"00",X"CC",X"CC",X"CC",X"00",X"00",X"00",X"0C",X"CC",X"C0",X"00",X"00",X"00",
		X"0C",X"CC",X"C0",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"0C",X"CC",X"C0",X"00",
		X"00",X"00",X"CC",X"CC",X"CC",X"00",X"00",X"0C",X"CC",X"CC",X"CC",X"C0",X"00",X"0C",X"CC",X"CC",
		X"CC",X"C0",X"00",X"0C",X"CC",X"CC",X"CC",X"C0",X"00",X"00",X"CC",X"CC",X"CC",X"00",X"00",X"00",
		X"0C",X"CC",X"C0",X"00",X"00",X"00",X"0C",X"00",X"C0",X"00",X"00",X"CC",X"CC",X"C0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"0C",X"CC",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",
		X"0C",X"CC",X"C0",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",
		X"00",X"00",X"0C",X"CC",X"C0",X"00",X"00",X"00",X"CC",X"CC",X"CC",X"00",X"00",X"00",X"CC",X"CC",
		X"CC",X"00",X"00",X"00",X"CC",X"CC",X"CC",X"00",X"00",X"00",X"0C",X"CC",X"C0",X"00",X"00",X"00",
		X"0C",X"0C",X"CC",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"CC",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"45",X"00",X"11",X"11",X"10",X"00",X"04",X"45",X"00",X"07",X"D1",
		X"00",X"00",X"05",X"54",X"45",X"EB",X"B7",X"00",X"00",X"00",X"55",X"44",X"AB",X"B7",X"00",X"00",
		X"00",X"0E",X"EE",X"AA",X"AA",X"A0",X"00",X"00",X"00",X"00",X"11",X"81",X"10",X"00",X"00",X"00",
		X"01",X"18",X"88",X"11",X"00",X"00",X"00",X"01",X"11",X"81",X"11",X"00",X"00",X"00",X"00",X"11",
		X"18",X"1A",X"00",X"00",X"00",X"01",X"18",X"81",X"11",X"00",X"00",X"00",X"01",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"11",X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",
		X"00",X"D1",X"1D",X"00",X"00",X"54",X"00",X"07",X"C0",X"00",X"00",X"E5",X"44",X"A7",X"70",X"00",
		X"00",X"0E",X"55",X"A7",X"71",X"10",X"00",X"00",X"01",X"16",X"81",X"10",X"00",X"00",X"00",X"16",
		X"11",X"00",X"00",X"00",X"01",X"11",X"61",X"10",X"00",X"00",X"01",X"11",X"11",X"10",X"00",X"00",
		X"00",X"10",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"11",X"00",X"54",X"50",X"00",X"00",
		X"1D",X"70",X"00",X"54",X"40",X"00",X"00",X"7B",X"BE",X"54",X"45",X"50",X"00",X"00",X"7B",X"BA",
		X"44",X"55",X"00",X"00",X"0A",X"AA",X"AA",X"EE",X"E0",X"00",X"00",X"01",X"18",X"11",X"00",X"00",
		X"00",X"00",X"11",X"88",X"81",X"10",X"00",X"00",X"00",X"11",X"18",X"11",X"10",X"00",X"00",X"00",
		X"A1",X"81",X"11",X"00",X"00",X"00",X"00",X"11",X"18",X"81",X"10",X"00",X"00",X"00",X"11",X"11",
		X"11",X"10",X"00",X"00",X"00",X"01",X"10",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0D",X"11",X"D0",X"04",X"40",X"00",X"00",X"C7",X"00",X"04",X"50",X"00",
		X"00",X"77",X"A4",X"45",X"E0",X"00",X"11",X"77",X"A5",X"5E",X"00",X"00",X"11",X"86",X"11",X"00",
		X"00",X"00",X"01",X"16",X"10",X"00",X"00",X"00",X"11",X"61",X"11",X"00",X"00",X"00",X"11",X"11",
		X"11",X"00",X"00",X"00",X"01",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",
		X"11",X"10",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"01",X"10",X"00",
		X"00",X"00",X"00",X"00",X"11",X"81",X"00",X"00",X"00",X"00",X"11",X"18",X"88",X"11",X"00",X"00",
		X"00",X"11",X"81",X"11",X"11",X"00",X"00",X"00",X"01",X"18",X"81",X"10",X"00",X"00",X"00",X"01",
		X"11",X"18",X"10",X"00",X"00",X"00",X"11",X"88",X"81",X"11",X"00",X"00",X"00",X"11",X"18",X"11",
		X"11",X"00",X"00",X"00",X"00",X"11",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"11",X"11",X"00",X"00",X"00",X"00",X"11",X"10",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"01",X"11",X"11",X"00",X"00",X"00",X"11",X"88",X"11",X"10",X"00",X"00",X"11",X"81",X"81",
		X"10",X"00",X"00",X"01",X"18",X"11",X"00",X"00",X"00",X"11",X"81",X"81",X"10",X"00",X"00",X"11",
		X"88",X"11",X"10",X"00",X"00",X"00",X"11",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"11",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"01",X"16",X"61",
		X"10",X"00",X"01",X"16",X"11",X"10",X"00",X"00",X"11",X"61",X"00",X"00",X"01",X"16",X"61",X"10",
		X"00",X"01",X"11",X"11",X"10",X"00",X"00",X"11",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"11",X"11",X"10",X"00",X"00",X"00",X"00",X"11",X"81",X"00",X"00",X"00",X"00",X"01",X"18",X"11",
		X"11",X"11",X"00",X"00",X"11",X"18",X"88",X"88",X"11",X"11",X"00",X"11",X"11",X"11",X"18",X"81",
		X"11",X"00",X"11",X"18",X"88",X"88",X"11",X"11",X"00",X"01",X"11",X"11",X"11",X"11",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"11",X"00",X"00",X"00",X"00",X"11",X"10",X"00",
		X"00",X"00",X"01",X"18",X"81",X"11",X"00",X"00",X"11",X"81",X"11",X"11",X"11",X"00",X"11",X"18",
		X"88",X"11",X"11",X"10",X"11",X"81",X"11",X"81",X"11",X"10",X"01",X"11",X"11",X"11",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"10",X"00",X"00",X"01",X"11",X"11",
		X"00",X"00",X"11",X"88",X"81",X"11",X"00",X"11",X"11",X"11",X"11",X"00",X"01",X"11",X"11",X"10",
		X"00",X"00",X"00",X"04",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"5E",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"68",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"E5",X"45",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5B",
		X"5E",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FA",X"AA",X"FF",X"70",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FD",X"47",X"77",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"05",
		X"22",X"4B",X"C7",X"7F",X"55",X"00",X"00",X"00",X"00",X"00",X"55",X"2F",X"E4",X"C7",X"F5",X"44",
		X"50",X"00",X"00",X"00",X"00",X"55",X"FF",X"77",X"FF",X"55",X"54",X"50",X"00",X"00",X"00",X"00",
		X"55",X"4B",X"FF",X"FB",X"4E",X"54",X"40",X"00",X"00",X"00",X"00",X"45",X"4B",X"BF",X"B4",X"2E",
		X"E5",X"45",X"00",X"00",X"00",X"00",X"45",X"EB",X"BF",X"B4",X"2E",X"EF",X"44",X"00",X"00",X"00",
		X"00",X"45",X"EF",X"BF",X"BF",X"EE",X"F5",X"44",X"04",X"00",X"00",X"00",X"44",X"EE",X"FF",X"F5",
		X"5E",X"54",X"44",X"E0",X"40",X"00",X"D0",X"DC",X"55",X"44",X"45",X"5E",X"D4",X"40",X"0E",X"04",
		X"00",X"04",X"40",X"55",X"54",X"45",X"E5",X"5C",X"EE",X"E0",X"E4",X"00",X"40",X"40",X"EE",X"54",
		X"44",X"55",X"55",X"E0",X"00",X"00",X"00",X"00",X"00",X"0E",X"E5",X"44",X"E5",X"4E",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"55",X"5E",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"E4",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"40",X"D0",X"00",X"0D",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"DD",X"00",X"0D",
		X"D4",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"40",X"00",X"B0",X"45",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"00",X"04",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"5E",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"88",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"E4",X"5E",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"45",X"EF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"AA",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D4",X"D7",X"77",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"24",X"47",X"77",X"F5",X"50",X"00",X"00",X"00",X"00",X"00",X"02",X"04",X"4E",
		X"7E",X"F4",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"BE",X"7F",X"54",X"44",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"7F",X"F5",X"55",X"44",X"50",X"00",X"00",X"00",X"00",X"00",X"00",
		X"54",X"25",X"5F",X"54",X"45",X"00",X"00",X"00",X"00",X"00",X"0E",X"B4",X"25",X"5F",X"54",X"45",
		X"00",X"00",X"00",X"00",X"0D",X"0E",X"B4",X"F5",X"5F",X"54",X"45",X"00",X"04",X"00",X"00",X"00",
		X"4E",X"BF",X"E5",X"F5",X"44",X"BE",X"E0",X"05",X"40",X"00",X"04",X"0E",X"FE",X"55",X"ED",X"4B",
		X"EE",X"EE",X"00",X"E0",X"00",X"00",X"05",X"E5",X"55",X"55",X"CE",X"EE",X"5E",X"0E",X"00",X"00",
		X"00",X"00",X"5E",X"5E",X"55",X"EE",X"E5",X"4E",X"E0",X"00",X"00",X"00",X"00",X"5E",X"EE",X"54",
		X"EE",X"54",X"EE",X"00",X"00",X"00",X"00",X"00",X"05",X"5E",X"5E",X"EE",X"EE",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"EE",X"45",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"B4",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"DD",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"B4",X"DD",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"44",X"00",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"04",X"50",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"5E",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"86",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"E5",X"55",X"4E",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"F5",X"54",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"AA",X"AF",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"D5",X"DD",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"77",X"75",X"42",X"2F",X"55",X"00",X"00",X"00",X"00",X"00",X"55",X"FF",X"75",X"4F",
		X"25",X"44",X"50",X"00",X"00",X"00",X"00",X"55",X"EF",X"F7",X"7F",X"55",X"54",X"50",X"00",X"00",
		X"00",X"00",X"55",X"4B",X"FF",X"FB",X"4E",X"54",X"40",X"00",X"00",X"00",X"00",X"45",X"4B",X"BF",
		X"B4",X"2E",X"E5",X"45",X"00",X"00",X"00",X"00",X"45",X"EB",X"BF",X"B4",X"2E",X"EF",X"44",X"00",
		X"00",X"00",X"00",X"45",X"EF",X"BF",X"BF",X"EE",X"F5",X"44",X"00",X"00",X"00",X"00",X"44",X"EE",
		X"FF",X"F5",X"5E",X"54",X"44",X"00",X"00",X"00",X"D0",X"DC",X"55",X"44",X"45",X"5E",X"D4",X"40",
		X"00",X"04",X"00",X"04",X"40",X"55",X"54",X"45",X"E5",X"5C",X"E0",X"0E",X"50",X"00",X"40",X"40",
		X"EE",X"54",X"44",X"55",X"55",X"EE",X"EE",X"04",X"00",X"00",X"00",X"0E",X"E5",X"44",X"E5",X"4E",
		X"E0",X"00",X"40",X"00",X"00",X"00",X"00",X"EE",X"55",X"5E",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"EE",X"E4",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"4D",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0D",X"D0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"B0",X"B4",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"45",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"5E",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"86",X"68",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"E5",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"54",X"45",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"7F",X"FF",X"EF",X"F7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"F2",X"4F",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"F7",X"02",X"2E",X"7F",X"40",X"00",X"00",X"00",X"00",
		X"00",X"5E",X"EE",X"50",X"5E",X"FE",X"54",X"00",X"00",X"00",X"00",X"05",X"5E",X"5F",X"F7",X"74",
		X"F5",X"E5",X"50",X"00",X"00",X"00",X"05",X"E5",X"4B",X"EF",X"FB",X"45",X"E5",X"40",X"00",X"00",
		X"00",X"05",X"E5",X"4B",X"BF",X"BB",X"E2",X"5E",X"45",X"00",X"00",X"00",X"04",X"E5",X"5B",X"BF",
		X"BB",X"52",X"5F",X"45",X"00",X"00",X"00",X"04",X"45",X"5F",X"BF",X"BF",X"55",X"5E",X"45",X"00",
		X"00",X"00",X"DE",X"CE",X"55",X"FF",X"F5",X"55",X"5E",X"40",X"00",X"00",X"00",X"0B",X"BE",X"E5",
		X"54",X"54",X"45",X"5D",X"00",X"00",X"00",X"00",X"B0",X"BE",X"E5",X"54",X"44",X"4E",X"5E",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"EE",X"55",X"44",X"E5",X"45",X"00",X"00",X"00",X"00",X"00",X"0E",
		X"EE",X"54",X"55",X"55",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"5E",X"EE",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4E",X"E4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0B",X"40",X"0B",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"0D",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"5D",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"45",X"04",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"44",X"B0",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E4",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"88",X"68",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"E5",X"45",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"EE",X"5B",X"50",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"7F",X"FA",X"AA",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"77",X"77",X"4D",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"05",X"5F",X"77",X"CB",X"42",X"25",X"00",X"00",X"00",X"00",X"00",
		X"54",X"45",X"F7",X"C4",X"EF",X"25",X"50",X"00",X"00",X"00",X"00",X"54",X"55",X"5F",X"F7",X"7F",
		X"F5",X"50",X"00",X"00",X"00",X"00",X"44",X"5E",X"4B",X"FF",X"FB",X"45",X"50",X"00",X"00",X"00",
		X"05",X"45",X"EE",X"24",X"BF",X"BB",X"45",X"40",X"00",X"00",X"00",X"04",X"4F",X"EE",X"24",X"BF",
		X"BB",X"E5",X"40",X"00",X"00",X"04",X"04",X"4E",X"EE",X"EF",X"BF",X"BF",X"E5",X"40",X"00",X"00",
		X"40",X"E4",X"4E",X"EE",X"55",X"FF",X"FE",X"E4",X"50",X"00",X"04",X"0E",X"D0",X"CE",X"EE",X"55",
		X"44",X"45",X"5D",X"00",X"00",X"04",X"E0",X"EB",X"BE",X"55",X"E5",X"44",X"55",X"55",X"00",X"00",
		X"00",X"00",X"B0",X"B5",X"55",X"54",X"44",X"55",X"45",X"00",X"00",X"00",X"00",X"00",X"EE",X"45",
		X"E4",X"45",X"E5",X"50",X"00",X"00",X"00",X"00",X"00",X"0E",X"EE",X"55",X"5E",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E4",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"B0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"0D",X"00",X"00",X"D0",X"4B",X"00",X"00",X"00",X"00",X"00",X"04",
		X"DD",X"00",X"0D",X"D4",X"40",X"00",X"00",X"00",X"00",X"00",X"05",X"40",X"B0",X"00",X"45",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E5",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"55",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"98",X"86",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"54",X"E5",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"E5",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F7",X"77",X"D4",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"F7",X"77",X"44",X"22",
		X"00",X"00",X"00",X"00",X"00",X"05",X"44",X"FE",X"7E",X"44",X"02",X"00",X"00",X"00",X"00",X"00",
		X"04",X"44",X"5F",X"7E",X"BE",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"45",X"55",X"FF",X"77",
		X"00",X"00",X"00",X"00",X"00",X"05",X"44",X"5F",X"55",X"24",X"50",X"00",X"00",X"00",X"00",X"00",
		X"05",X"44",X"5F",X"55",X"24",X"BE",X"00",X"00",X"00",X"04",X"00",X"05",X"44",X"5F",X"55",X"F4",
		X"BE",X"00",X"00",X"00",X"45",X"00",X"EE",X"D4",X"CE",X"E5",X"EF",X"BE",X"00",X"00",X"00",X"E0",
		X"0E",X"EE",X"EB",X"BE",X"E5",X"5E",X"FE",X"00",X"00",X"00",X"0E",X"0E",X"5E",X"BE",X"B5",X"55",
		X"55",X"E5",X"00",X"00",X"00",X"00",X"EE",X"45",X"EE",X"E5",X"5E",X"5E",X"50",X"00",X"00",X"00",
		X"00",X"0E",X"E4",X"5E",X"E4",X"5E",X"EE",X"50",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",
		X"5E",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"E5",X"4E",X"E5",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0D",X"04",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4D",X"D0",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"D0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"40",X"0D",X"D4",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",
		X"04",X"44",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"54",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"55",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"86",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"45",X"55",
		X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E4",X"55",X"FF",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"AA",X"AF",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"D5",
		X"D7",X"70",X"00",X"00",X"00",X"00",X"00",X"05",X"5F",X"22",X"45",X"77",X"75",X"00",X"00",X"00",
		X"00",X"00",X"54",X"45",X"2F",X"45",X"7F",X"F5",X"50",X"00",X"00",X"00",X"00",X"54",X"55",X"5F",
		X"77",X"FF",X"E5",X"50",X"00",X"00",X"00",X"00",X"44",X"5E",X"4B",X"FF",X"FB",X"45",X"50",X"00",
		X"00",X"00",X"05",X"45",X"EE",X"24",X"BF",X"BB",X"45",X"40",X"00",X"00",X"00",X"04",X"4F",X"EE",
		X"24",X"BF",X"BB",X"E5",X"40",X"00",X"00",X"00",X"04",X"4E",X"EE",X"EF",X"BF",X"BF",X"E5",X"40",
		X"00",X"00",X"00",X"04",X"4E",X"EE",X"55",X"FF",X"FE",X"E4",X"50",X"00",X"04",X"00",X"DF",X"CE",
		X"EE",X"55",X"44",X"45",X"5D",X"00",X"00",X"00",X"5E",X"0B",X"BE",X"55",X"E5",X"44",X"55",X"55",
		X"00",X"00",X"04",X"0E",X"BE",X"BE",X"55",X"54",X"44",X"55",X"45",X"00",X"00",X"00",X"40",X"00",
		X"EE",X"45",X"E4",X"45",X"E5",X"50",X"00",X"00",X"00",X"00",X"00",X"0E",X"EE",X"55",X"5E",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E4",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"4B",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"4D",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"44",X"B0",X"B0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"50",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",
		X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"08",X"66",X"80",X"50",X"00",X"00",
		X"00",X"00",X"05",X"55",X"5F",X"55",X"55",X"5E",X"00",X"55",X"00",X"00",X"00",X"54",X"44",X"5F",
		X"F5",X"44",X"5F",X"F4",X"44",X"50",X"00",X"05",X"44",X"04",X"F7",X"FF",X"FE",X"FF",X"7E",X"04",
		X"45",X"00",X"04",X"40",X"55",X"E7",X"7F",X"25",X"F7",X"7E",X"50",X"44",X"00",X"04",X"45",X"55",
		X"5E",X"7F",X"22",X"07",X"E5",X"55",X"44",X"00",X"DE",X"CE",X"55",X"EE",X"FF",X"FF",X"F0",X"E5",
		X"5E",X"CE",X"00",X"0B",X"BE",X"E5",X"E4",X"BB",X"FB",X"B4",X"25",X"EE",X"BB",X"00",X"B0",X"BE",
		X"E5",X"5E",X"BB",X"FB",X"BE",X"2E",X"EB",X"EB",X"B0",X"00",X"EE",X"55",X"55",X"FB",X"FB",X"F5",
		X"55",X"EE",X"E0",X"00",X"00",X"EE",X"55",X"54",X"4F",X"FF",X"54",X"45",X"5E",X"00",X"00",X"00",
		X"0E",X"E5",X"54",X"45",X"55",X"54",X"45",X"5E",X"00",X"00",X"00",X"0E",X"EE",X"55",X"44",X"55",
		X"44",X"5E",X"E0",X"00",X"00",X"00",X"00",X"EE",X"EE",X"55",X"45",X"55",X"EE",X"E0",X"00",X"00",
		X"00",X"00",X"0E",X"EE",X"EE",X"EE",X"EE",X"E0",X"00",X"00",X"00",X"00",X"40",X"00",X"B4",X"4E",
		X"EE",X"44",X"B0",X"00",X"40",X"00",X"00",X"44",X"0D",X"40",X"00",X"00",X"00",X"4D",X"04",X"40",
		X"00",X"00",X"04",X"DD",X"00",X"00",X"00",X"00",X"0D",X"D4",X"00",X"00",X"00",X"44",X"40",X"00",
		X"00",X"00",X"00",X"00",X"44",X"40",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"05",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",
		X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"54",X"EE",X"EE",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"45",X"AA",X"F7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F2",X"47",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"27",X"4E",X"7F",X"55",X"50",X"00",X"00",X"00",X"00",
		X"55",X"FF",X"47",X"F5",X"E4",X"45",X"00",X"00",X"00",X"00",X"55",X"44",X"FF",X"4E",X"E5",X"45",
		X"00",X"00",X"00",X"00",X"55",X"BB",X"FB",X"42",X"5E",X"44",X"50",X"00",X"00",X"00",X"4E",X"BB",
		X"FB",X"B5",X"5E",X"E4",X"50",X"00",X"00",X"00",X"4E",X"FB",X"FB",X"F5",X"5E",X"F4",X"40",X"00",
		X"00",X"00",X"4E",X"EF",X"FF",X"55",X"5E",X"44",X"40",X"40",X"00",X"D0",X"D5",X"E5",X"44",X"55",
		X"ED",X"44",X"E0",X"04",X"00",X"04",X"40",X"E5",X"44",X"5E",X"55",X"C0",X"0E",X"04",X"00",X"05",
		X"50",X"EE",X"54",X"4F",X"55",X"5E",X"EE",X"04",X"00",X"00",X"00",X"0E",X"E5",X"5F",X"54",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"55",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"E4",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"D4",X"04",X"00",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"E4",X"D0",X"00",X"D4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"5E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5E",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"4F",X"FF",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"77",X"70",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"D4",X"E7",X"75",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E4",X"E7",X"F5",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"F5",X"E5",X"44",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"B5",X"5E",X"54",X"40",X"00",X"00",X"00",X"00",X"00",X"EB",X"42",
		X"5E",X"55",X"45",X"00",X"00",X"00",X"00",X"D0",X"EB",X"45",X"55",X"E4",X"45",X"00",X"00",X"00",
		X"00",X"04",X"E4",X"F5",X"55",X"44",X"4E",X"00",X"05",X"00",X"00",X"05",X"5F",X"55",X"5E",X"D4",
		X"55",X"E0",X"05",X"40",X"00",X"00",X"0E",X"55",X"E5",X"5C",X"FE",X"EE",X"0E",X"00",X"00",X"00",
		X"05",X"EE",X"F5",X"4F",X"E5",X"5E",X"E0",X"00",X"00",X"00",X"00",X"5E",X"EF",X"EE",X"E5",X"4E",
		X"00",X"00",X"00",X"00",X"00",X"05",X"5E",X"EE",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"E4",X"E0",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"5D",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"4D",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"44",
		X"40",X"04",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"5E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"86",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"E5",X"54",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7A",
		X"AE",X"5A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"F2",X"FA",X"50",X"00",X"00",X"00",
		X"00",X"00",X"05",X"F7",X"4E",X"2F",X"55",X"50",X"00",X"00",X"00",X"00",X"55",X"5F",X"47",X"F5",
		X"E4",X"45",X"00",X"00",X"00",X"00",X"55",X"44",X"FF",X"4E",X"E5",X"45",X"00",X"00",X"00",X"00",
		X"55",X"BB",X"FB",X"42",X"5E",X"44",X"50",X"00",X"00",X"00",X"4E",X"BB",X"FB",X"B5",X"5E",X"E4",
		X"50",X"00",X"00",X"00",X"4E",X"FB",X"FB",X"F5",X"5E",X"F4",X"40",X"00",X"00",X"00",X"4E",X"EF",
		X"FF",X"55",X"5E",X"44",X"40",X"00",X"00",X"D0",X"D5",X"E5",X"44",X"55",X"ED",X"44",X"E0",X"00",
		X"00",X"04",X"40",X"E5",X"44",X"5E",X"55",X"C0",X"00",X"00",X"00",X"05",X"50",X"EE",X"54",X"4F",
		X"55",X"5E",X"E0",X"50",X"00",X"00",X"00",X"0E",X"E5",X"5F",X"54",X"E0",X"0E",X"04",X"00",X"00",
		X"00",X"00",X"EE",X"55",X"EE",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"0E",X"E4",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0D",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4D",X"50",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"04",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"5E",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"86",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E5",X"55",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"79",X"A4",X"5A",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"92",X"4F",X"70",X"00",X"00",
		X"00",X"00",X"00",X"05",X"F7",X"EE",X"57",X"FE",X"50",X"00",X"00",X"00",X"00",X"05",X"EF",X"E7",
		X"4F",X"EE",X"40",X"00",X"00",X"00",X"00",X"EE",X"44",X"FF",X"F4",X"45",X"55",X"00",X"00",X"00",
		X"00",X"5E",X"4B",X"BF",X"B4",X"42",X"E4",X"00",X"00",X"00",X"00",X"4E",X"EB",X"BF",X"BB",X"55",
		X"EE",X"50",X"00",X"00",X"00",X"4E",X"EF",X"BF",X"BF",X"55",X"5E",X"50",X"00",X"00",X"00",X"4E",
		X"E5",X"FF",X"F5",X"55",X"5E",X"40",X"00",X"00",X"D0",X"D5",X"E5",X"44",X"44",X"55",X"5D",X"40",
		X"00",X"00",X"04",X"4E",X"E5",X"54",X"44",X"5E",X"55",X"00",X"00",X"00",X"0E",X"EE",X"EE",X"54",
		X"45",X"5E",X"54",X"00",X"00",X"00",X"00",X"00",X"EE",X"E5",X"5E",X"EE",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"EE",X"5E",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4E",X"E4",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"D0",X"0D",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"45",X"54",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"E5",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"86",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"EE",X"E4",X"5E",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"FA",X"A5",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"77",X"42",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"55",X"5F",X"7E",X"47",X"25",X"00",X"00",X"00",X"00",X"05",X"44",X"E5",X"F7",X"4F",X"F5",X"50",
		X"00",X"00",X"00",X"05",X"45",X"EE",X"4F",X"F4",X"45",X"50",X"00",X"00",X"00",X"54",X"4E",X"55",
		X"4B",X"FB",X"B2",X"50",X"00",X"00",X"00",X"54",X"EE",X"55",X"BB",X"FB",X"BE",X"40",X"00",X"00",
		X"00",X"44",X"FE",X"55",X"FB",X"FB",X"FE",X"40",X"00",X"00",X"40",X"44",X"EE",X"55",X"5F",X"FF",
		X"EE",X"40",X"00",X"04",X"0D",X"FC",X"E5",X"55",X"54",X"45",X"ED",X"00",X"00",X"04",X"0E",X"44",
		X"E5",X"55",X"54",X"45",X"E5",X"00",X"00",X"04",X"0E",X"55",X"EE",X"55",X"44",X"5E",X"45",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"55",X"55",X"EE",X"50",X"00",X"00",X"00",X"00",X"00",X"0E",X"E5",
		X"5E",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E4",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E0",X"04",X"04",X"D0",X"40",X"00",X"00",X"00",X"00",X"00",X"04",X"D0",X"00",X"D4",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"40",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"86",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"EE",X"EE",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",
		X"FF",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"77",X"74",X"20",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"44",X"77",X"E4",X"D2",X"00",X"00",X"00",X"00",X"00",X"04",X"44",X"F7",X"E4",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"54",X"45",X"E5",X"FF",X"70",X"00",X"00",X"00",X"00",X"00",X"44",
		X"EE",X"55",X"B5",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"EE",X"55",X"4B",X"E0",X"00",X"00",
		X"00",X"00",X"0E",X"44",X"E5",X"55",X"4B",X"E0",X"00",X"00",X"05",X"00",X"ED",X"FC",X"E5",X"55",
		X"F4",X"E0",X"00",X"00",X"45",X"0E",X"EE",X"BB",X"5E",X"55",X"5F",X"E0",X"00",X"00",X"0E",X"0E",
		X"5E",X"EE",X"E5",X"55",X"5E",X"00",X"00",X"00",X"00",X"EE",X"5E",X"E5",X"55",X"55",X"E5",X"00",
		X"00",X"00",X"00",X"0E",X"E5",X"EE",X"55",X"EE",X"50",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",
		X"EE",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"E4",X"E5",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"4D",X"5D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"0D",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"44",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"55",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",
		X"E4",X"55",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"5E",X"AA",X"70",X"00",X"00",X"00",
		X"00",X"00",X"00",X"5A",X"F2",X"F7",X"70",X"00",X"00",X"00",X"00",X"00",X"55",X"5F",X"2E",X"47",
		X"F5",X"00",X"00",X"00",X"00",X"05",X"44",X"E5",X"F7",X"4F",X"55",X"50",X"00",X"00",X"00",X"05",
		X"45",X"EE",X"4F",X"F4",X"45",X"50",X"00",X"00",X"00",X"54",X"4E",X"55",X"4B",X"FB",X"B2",X"50",
		X"00",X"00",X"00",X"54",X"EE",X"55",X"BB",X"FB",X"BE",X"40",X"00",X"00",X"00",X"44",X"FE",X"55",
		X"FB",X"FB",X"FE",X"40",X"00",X"00",X"00",X"44",X"EE",X"55",X"5F",X"FF",X"EE",X"40",X"00",X"00",
		X"0D",X"FC",X"E5",X"55",X"54",X"45",X"ED",X"00",X"00",X"00",X"00",X"44",X"E5",X"55",X"54",X"45",
		X"E5",X"00",X"00",X"00",X"50",X"55",X"EE",X"55",X"44",X"5E",X"45",X"00",X"00",X"04",X"0E",X"00",
		X"EE",X"55",X"55",X"EE",X"50",X"00",X"00",X"00",X"50",X"00",X"0E",X"E5",X"5E",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E4",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4D",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"5D",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"68",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"55",X"5E",X"EE",X"00",X"00",X"00",X"00",X"05",X"45",X"07",X"AA",
		X"45",X"A7",X"45",X"00",X"00",X"00",X"54",X"4E",X"F7",X"7A",X"24",X"F7",X"F4",X"50",X"00",X"05",
		X"45",X"55",X"EF",X"7E",X"E5",X"7F",X"EE",X"45",X"00",X"05",X"4E",X"54",X"44",X"FE",X"74",X"F4",
		X"2E",X"44",X"00",X"05",X"4E",X"54",X"4B",X"BF",X"FF",X"BB",X"4F",X"44",X"00",X"D0",X"DE",X"55",
		X"FB",X"BB",X"FB",X"BB",X"FB",X"DD",X"00",X"0B",X"BE",X"E5",X"5F",X"BB",X"FB",X"BF",X"5B",X"EB",
		X"00",X"00",X"0E",X"E5",X"55",X"5F",X"FF",X"55",X"5E",X"E0",X"00",X"00",X"00",X"EE",X"55",X"54",
		X"44",X"55",X"EE",X"00",X"00",X"00",X"00",X"0E",X"E5",X"55",X"45",X"EE",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"EE",X"EE",X"E0",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"00",X"04",
		X"00",X"04",X"00",X"00",X"04",X"D4",X"00",X"00",X"00",X"00",X"4D",X"40",X"00",X"00",X"44",X"4D",
		X"00",X"00",X"00",X"00",X"D4",X"44",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"5E",X"EF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"68",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"F5",X"45",X"5E",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"AA",X"A7",X"F0",X"00",X"00",X"00",X"00",X"00",X"F2",X"D7",
		X"77",X"FF",X"00",X"00",X"00",X"00",X"0F",X"52",X"F4",X"7F",X"55",X"F0",X"00",X"00",X"00",X"FE",
		X"5F",X"FF",X"FE",X"54",X"5F",X"00",X"00",X"00",X"F5",X"BB",X"FB",X"B2",X"E4",X"4F",X"00",X"00",
		X"00",X"F5",X"4B",X"FB",X"45",X"EF",X"45",X"F0",X"00",X"00",X"F5",X"EF",X"BF",X"E5",X"EF",X"45",
		X"F0",X"00",X"00",X"F4",X"EE",X"F5",X"55",X"54",X"4F",X"4F",X"00",X"00",X"D7",X"EE",X"54",X"55",
		X"D4",X"5F",X"F4",X"F0",X"00",X"E7",X"EE",X"54",X"5F",X"5C",X"EE",X"E4",X"F0",X"00",X"FF",X"FE",
		X"E5",X"5F",X"45",X"EF",X"FF",X"00",X"00",X"00",X"0F",X"EE",X"5E",X"FE",X"EF",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"EE",X"5E",X"F0",X"00",X"00",X"00",X"00",X"0F",X"50",X"F5",X"F4",X"FF",X"00",
		X"00",X"00",X"00",X"0F",X"45",X"DF",X"0F",X"D5",X"F0",X"00",X"00",X"00",X"00",X"F4",X"5F",X"00",
		X"F4",X"F0",X"00",X"00",X"00",X"00",X"0F",X"F4",X"FF",X"45",X"F0",X"00",X"00",X"00",X"FF",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"55",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"68",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"F5",X"EE",X"EE",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"FF",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"F2",X"24",X"77",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"F2",X"F4",X"57",X"55",X"F0",X"00",X"00",X"00",X"00",X"0F",X"77",X"FE",X"54",
		X"5F",X"00",X"00",X"00",X"00",X"00",X"FF",X"5E",X"E4",X"45",X"F0",X"00",X"00",X"00",X"0F",X"EB",
		X"25",X"EE",X"44",X"F0",X"00",X"00",X"00",X"D4",X"BB",X"55",X"EE",X"44",X"F0",X"00",X"00",X"00",
		X"F5",X"B5",X"55",X"E4",X"45",X"F0",X"0F",X"00",X"00",X"0F",X"5E",X"5E",X"5D",X"CE",X"EF",X"F5",
		X"F0",X"00",X"0F",X"FE",X"EE",X"55",X"EE",X"5E",X"F5",X"40",X"00",X"00",X"F5",X"EE",X"45",X"E5",
		X"5E",X"FE",X"F0",X"00",X"00",X"0F",X"5E",X"EE",X"EE",X"EE",X"EF",X"00",X"00",X"00",X"00",X"FF",
		X"5E",X"4E",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"4F",X"D4",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"F4",X"D0",X"F4",X"F0",X"00",X"00",X"00",X"00",X"0F",X"4F",X"44",X"FF",X"40",X"00",
		X"00",X"00",X"0F",X"5E",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"58",X"6F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F5",X"55",X"4E",X"F0",X"00",X"00",X"00",X"00",X"00",X"07",X"AA",X"AF",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"F7",X"74",X"22",X"FF",X"00",X"00",X"00",X"00",X"0F",X"5F",
		X"74",X"52",X"55",X"F0",X"00",X"00",X"00",X"FE",X"5F",X"FF",X"FE",X"54",X"5F",X"00",X"00",X"00",
		X"F5",X"BB",X"FB",X"B2",X"E4",X"4F",X"00",X"00",X"00",X"F5",X"4B",X"FB",X"45",X"EF",X"45",X"F0",
		X"00",X"00",X"F5",X"EF",X"BF",X"E5",X"EF",X"45",X"F0",X"00",X"00",X"F4",X"EE",X"F5",X"55",X"54",
		X"4F",X"00",X"00",X"00",X"D7",X"EE",X"54",X"55",X"D4",X"5F",X"F0",X"F0",X"00",X"E7",X"EE",X"54",
		X"5F",X"5C",X"EE",X"EF",X"50",X"00",X"FF",X"FE",X"E5",X"5F",X"45",X"EF",X"F4",X"F0",X"00",X"00",
		X"0F",X"EE",X"5E",X"FE",X"EF",X"0F",X"00",X"00",X"00",X"00",X"FE",X"EE",X"5E",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"F4",X"4F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"D4",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F4",X"DF",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"4F",
		X"44",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"5E",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"86",X"EF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F5",X"54",X"5E",X"00",X"00",X"00",X"00",X"00",X"00",X"FA",X"AA",X"AA",X"F0",X"00",
		X"00",X"00",X"00",X"0F",X"F7",X"E2",X"E7",X"FF",X"00",X"00",X"00",X"00",X"FE",X"E7",X"72",X"47",
		X"55",X"F0",X"00",X"00",X"0F",X"EE",X"EE",X"F7",X"F5",X"E5",X"5F",X"00",X"00",X"0F",X"5E",X"E4",
		X"BE",X"4B",X"2E",X"5F",X"00",X"00",X"0F",X"5E",X"E4",X"BF",X"4B",X"EE",X"5F",X"00",X"00",X"0F",
		X"5E",X"EE",X"FB",X"F5",X"EE",X"4F",X"00",X"00",X"0F",X"4E",X"EE",X"5F",X"55",X"5E",X"4F",X"00",
		X"00",X"0D",X"7E",X"5E",X"55",X"45",X"5E",X"DF",X"00",X"00",X"0F",X"7E",X"E5",X"55",X"45",X"55",
		X"EF",X"00",X"00",X"00",X"FF",X"EE",X"E5",X"55",X"E5",X"EF",X"00",X"00",X"00",X"00",X"FE",X"E5",
		X"5E",X"EE",X"F0",X"00",X"00",X"00",X"00",X"0F",X"EE",X"EE",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"4F",X"F4",X"F0",X"00",X"00",X"00",X"00",X"00",X"F5",X"DF",X"FD",X"5F",X"00",X"00",X"00",
		X"00",X"0F",X"44",X"F4",X"4F",X"44",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"E5",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"86",X"F0",X"00",X"00",X"00",X"00",X"00",X"0F",X"E5",
		X"54",X"5F",X"00",X"00",X"00",X"00",X"00",X"0F",X"7A",X"AA",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"77",X"7D",X"2F",X"00",X"00",X"00",X"00",X"0F",X"55",X"F7",X"4F",X"25",X"F0",X"00",X"00",
		X"00",X"F5",X"45",X"EF",X"FF",X"F5",X"EF",X"00",X"00",X"00",X"F4",X"4E",X"5B",X"BF",X"B2",X"5F",
		X"00",X"00",X"0F",X"54",X"FE",X"54",X"BF",X"B4",X"5F",X"00",X"00",X"0F",X"54",X"FE",X"5E",X"FB",
		X"FE",X"5F",X"00",X"00",X"F4",X"F4",X"45",X"55",X"5F",X"EE",X"4F",X"00",X"0F",X"4F",X"FD",X"7E",
		X"55",X"45",X"EE",X"4F",X"00",X"0F",X"4E",X"EE",X"75",X"E5",X"45",X"E5",X"F0",X"00",X"00",X"FF",
		X"FE",X"5E",X"E5",X"5E",X"E5",X"F0",X"00",X"00",X"00",X"FE",X"EE",X"E5",X"EE",X"FF",X"00",X"00",
		X"00",X"00",X"0F",X"E5",X"EE",X"EF",X"00",X"00",X"00",X"00",X"00",X"FF",X"4F",X"5F",X"05",X"F0",
		X"00",X"00",X"00",X"0F",X"5D",X"F0",X"FD",X"54",X"F0",X"00",X"00",X"00",X"0F",X"4F",X"00",X"F5",
		X"4F",X"00",X"00",X"00",X"00",X"0F",X"54",X"FF",X"4F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"55",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FE",X"86",X"F0",X"00",X"00",X"00",X"00",X"00",X"0F",X"EE",X"EE",X"5F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"FF",X"77",
		X"42",X"2F",X"00",X"00",X"00",X"00",X"0F",X"55",X"75",X"4F",X"2F",X"00",X"00",X"00",X"00",X"F5",
		X"45",X"EF",X"77",X"F0",X"00",X"00",X"00",X"0F",X"54",X"4E",X"E5",X"FF",X"00",X"00",X"00",X"00",
		X"0F",X"44",X"EE",X"55",X"BE",X"F0",X"00",X"00",X"00",X"0F",X"44",X"EE",X"55",X"BB",X"F0",X"00",
		X"00",X"F0",X"0F",X"D7",X"EE",X"55",X"5B",X"F0",X"00",X"0F",X"5F",X"FE",X"E7",X"E5",X"E5",X"E5",
		X"F0",X"00",X"04",X"5F",X"E5",X"EE",X"55",X"EE",X"EF",X"F0",X"00",X"0F",X"EF",X"E5",X"5E",X"54",
		X"EE",X"5F",X"00",X"00",X"00",X"FE",X"EE",X"EE",X"EE",X"E5",X"F0",X"00",X"00",X"00",X"00",X"FE",
		X"E4",X"E5",X"FF",X"00",X"00",X"00",X"00",X"0F",X"4D",X"F4",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"4F",X"0D",X"4F",X"00",X"00",X"00",X"00",X"00",X"04",X"FF",X"44",X"F4",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FE",X"E5",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"F6",X"8E",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"0F",X"E4",X"5E",X"EF",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"FA",X"AA",X"70",X"00",X"00",X"00",X"00",X"00",X"FF",X"22",X"47",X"7F",X"00",X"00",X"00",X"00",
		X"0F",X"55",X"25",X"47",X"F5",X"F0",X"00",X"00",X"00",X"F5",X"45",X"EF",X"FF",X"F5",X"EF",X"00",
		X"00",X"00",X"F4",X"4E",X"5B",X"BF",X"B2",X"5F",X"00",X"00",X"0F",X"54",X"FE",X"54",X"BF",X"B4",
		X"5F",X"00",X"00",X"0F",X"54",X"FE",X"5E",X"FB",X"FE",X"5F",X"00",X"00",X"00",X"F4",X"45",X"55",
		X"5F",X"EE",X"4F",X"00",X"0F",X"0F",X"FD",X"7E",X"55",X"45",X"EE",X"4F",X"00",X"05",X"FE",X"EE",
		X"75",X"E5",X"45",X"E5",X"F0",X"00",X"0F",X"4F",X"FE",X"5E",X"E5",X"5E",X"E5",X"F0",X"00",X"00",
		X"F0",X"FE",X"EE",X"E5",X"EE",X"F0",X"00",X"00",X"00",X"00",X"0F",X"E5",X"EE",X"EF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F4",X"4F",X"F0",X"00",X"00",X"00",X"00",X"00",X"0F",X"4D",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"4F",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"44",
		X"F4",X"F0",X"00",X"00",X"00",X"00",X"00",X"0F",X"5E",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"86",X"EF",X"00",X"00",X"00",X"00",X"00",X"0F",X"F5",X"54",X"5E",X"FF",X"00",X"00",X"00",
		X"0F",X"F5",X"09",X"99",X"99",X"05",X"FF",X"00",X"00",X"F5",X"45",X"E7",X"E2",X"E7",X"E5",X"45",
		X"F0",X"00",X"54",X"EE",X"E7",X"72",X"47",X"EE",X"E4",X"5F",X"00",X"54",X"4E",X"EE",X"F0",X"FE",
		X"2E",X"44",X"5F",X"00",X"D7",X"E5",X"E4",X"BF",X"4B",X"E5",X"ED",X"7F",X"00",X"F7",X"55",X"EE",
		X"BF",X"BE",X"E5",X"7E",X"7F",X"00",X"FE",X"E5",X"55",X"5F",X"55",X"55",X"EE",X"F0",X"00",X"0F",
		X"EE",X"55",X"55",X"55",X"5E",X"EF",X"00",X"00",X"00",X"FF",X"EE",X"EE",X"EE",X"EF",X"F0",X"00",
		X"00",X"F4",X"0F",X"4F",X"FF",X"FF",X"4F",X"04",X"F0",X"00",X"0F",X"4D",X"F0",X"00",X"00",X"FD",
		X"4F",X"00",X"00",X"0F",X"4F",X"00",X"00",X"00",X"0F",X"4F",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"0E",X"EE",X"E0",X"BB",
		X"B0",X"00",X"00",X"05",X"05",X"00",X"05",X"00",X"DD",X"D0",X"00",X"00",X"04",X"00",X"0E",X"4E",
		X"40",X"33",X"30",X"00",X"00",X"BB",X"B0",X"EE",X"EE",X"00",X"E0",X"00",X"00",X"00",X"DD",X"D0",
		X"05",X"00",X"05",X"05",X"00",X"00",X"00",X"33",X"30",X"4E",X"4E",X"00",X"04",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"00",X"09",X"99",X"9A",X"00",X"00",X"00",X"00",X"9A",X"A0",X"00",X"00",
		X"00",X"09",X"88",X"90",X"00",X"00",X"00",X"00",X"88",X"9A",X"00",X"00",X"00",X"00",X"00",X"89",
		X"A0",X"00",X"00",X"00",X"0C",X"99",X"9A",X"00",X"00",X"00",X"0E",X"99",X"A9",X"A0",X"00",X"00",
		X"09",X"9A",X"0A",X"90",X"00",X"00",X"A9",X"9A",X"09",X"90",X"00",X"09",X"A9",X"9A",X"88",X"00",
		X"00",X"89",X"09",X"9A",X"A0",X"00",X"00",X"00",X"00",X"A8",X"99",X"00",X"00",X"00",X"00",X"98",
		X"99",X"00",X"00",X"00",X"09",X"9A",X"00",X"00",X"00",X"90",X"99",X"A0",X"A9",X"A0",X"00",X"A9",
		X"90",X"00",X"00",X"99",X"00",X"00",X"90",X"00",X"09",X"90",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"09",X"99",X"9A",X"00",X"00",X"00",X"00",X"9A",X"A0",X"00",X"00",X"00",X"09",X"88",X"90",
		X"00",X"00",X"00",X"00",X"88",X"9A",X"00",X"00",X"00",X"00",X"00",X"89",X"00",X"00",X"00",X"00",
		X"0C",X"99",X"A0",X"00",X"00",X"00",X"0E",X"99",X"90",X"00",X"00",X"00",X"09",X"9A",X"9A",X"00",
		X"00",X"00",X"09",X"9A",X"9A",X"00",X"00",X"00",X"09",X"99",X"90",X"00",X"00",X"00",X"09",X"98",
		X"80",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"89",X"90",X"00",X"00",X"00",
		X"00",X"89",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A9",X"00",X"00",
		X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"09",X"99",X"9A",
		X"00",X"00",X"00",X"00",X"9A",X"A0",X"00",X"00",X"00",X"09",X"88",X"90",X"00",X"00",X"00",X"00",
		X"88",X"9A",X"00",X"00",X"00",X"00",X"00",X"89",X"00",X"00",X"00",X"00",X"0C",X"99",X"A0",X"00",
		X"00",X"00",X"0E",X"99",X"9A",X"00",X"00",X"00",X"09",X"90",X"09",X"00",X"00",X"00",X"09",X"9A",
		X"9A",X"00",X"00",X"00",X"09",X"88",X"90",X"00",X"00",X"00",X"09",X"A9",X"00",X"00",X"00",X"00",
		X"08",X"99",X"00",X"00",X"00",X"00",X"08",X"99",X"00",X"00",X"00",X"00",X"00",X"A9",X"90",X"00",
		X"00",X"00",X"0A",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"0A",X"9A",X"00",X"00",X"99",X"00",
		X"09",X"90",X"00",X"00",X"00",X"A9",X"A0",X"00",X"00",X"00",X"09",X"99",X"99",X"00",X"00",X"00",
		X"00",X"AA",X"A0",X"00",X"00",X"00",X"00",X"89",X"80",X"00",X"00",X"00",X"00",X"98",X"90",X"00",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"A9",X"8E",X"89",X"A0",X"00",X"00",X"99",X"9C",
		X"99",X"90",X"00",X"00",X"9A",X"99",X"9A",X"90",X"00",X"00",X"90",X"9A",X"90",X"90",X"00",X"00",
		X"90",X"9A",X"90",X"90",X"00",X"00",X"80",X"9A",X"90",X"80",X"00",X"00",X"00",X"0A",X"00",X"A0",
		X"00",X"00",X"00",X"09",X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"90",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"A9",X"A0",X"00",X"00",X"00",X"00",X"9A",X"90",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"A9",X"99",X"90",X"00",X"00",X"00",X"0A",X"A9",X"00",
		X"00",X"00",X"00",X"09",X"88",X"90",X"00",X"00",X"00",X"A9",X"88",X"00",X"00",X"00",X"0A",X"98",
		X"00",X"00",X"00",X"00",X"A9",X"99",X"C0",X"00",X"00",X"0A",X"9A",X"99",X"E0",X"00",X"00",X"09",
		X"A0",X"A9",X"90",X"00",X"00",X"09",X"90",X"A9",X"9A",X"00",X"00",X"00",X"88",X"A9",X"9A",X"90",
		X"00",X"00",X"0A",X"A9",X"90",X"98",X"00",X"00",X"99",X"8A",X"00",X"00",X"00",X"00",X"99",X"89",
		X"00",X"00",X"00",X"00",X"00",X"A9",X"90",X"00",X"00",X"0A",X"9A",X"0A",X"99",X"09",X"00",X"99",
		X"00",X"00",X"09",X"9A",X"00",X"09",X"90",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"A9",X"99",X"90",X"00",X"00",X"00",X"0A",X"A9",X"00",X"00",X"00",X"00",X"09",
		X"88",X"90",X"00",X"00",X"00",X"A9",X"88",X"00",X"00",X"00",X"00",X"98",X"00",X"00",X"00",X"00",
		X"0A",X"99",X"C0",X"00",X"00",X"00",X"09",X"99",X"E0",X"00",X"00",X"00",X"A9",X"A9",X"90",X"00",
		X"00",X"00",X"A9",X"A9",X"90",X"00",X"00",X"00",X"09",X"99",X"90",X"00",X"00",X"00",X"08",X"89",
		X"90",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"09",X"98",X"00",X"00",X"00",X"00",
		X"09",X"98",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9A",X"00",X"00",
		X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"A9",
		X"99",X"90",X"00",X"00",X"00",X"0A",X"A9",X"00",X"00",X"00",X"00",X"09",X"88",X"90",X"00",X"00",
		X"00",X"A9",X"88",X"00",X"00",X"00",X"00",X"98",X"00",X"00",X"00",X"00",X"0A",X"99",X"C0",X"00",
		X"00",X"00",X"A9",X"99",X"E0",X"00",X"00",X"00",X"90",X"09",X"90",X"00",X"00",X"00",X"A9",X"A9",
		X"90",X"00",X"00",X"00",X"09",X"88",X"90",X"00",X"00",X"00",X"00",X"9A",X"90",X"00",X"00",X"00",
		X"00",X"99",X"80",X"00",X"00",X"00",X"00",X"99",X"80",X"00",X"00",X"00",X"09",X"9A",X"00",X"00",
		X"00",X"00",X"99",X"00",X"A0",X"00",X"00",X"A9",X"A0",X"00",X"90",X"00",X"00",X"09",X"90",X"00",
		X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"A9",X"A0",X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"89",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"98",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"A9",X"E5",X"E9",X"A0",X"00",X"00",X"00",X"00",X"99",X"55",X"59",
		X"90",X"00",X"00",X"00",X"00",X"9A",X"55",X"5A",X"90",X"00",X"00",X"00",X"00",X"90",X"E5",X"E0",
		X"90",X"00",X"00",X"00",X"00",X"90",X"9E",X"90",X"90",X"00",X"00",X"00",X"00",X"80",X"9A",X"90",
		X"80",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"90",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"A9",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"9A",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"A9",X"A0",X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E5",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"94",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"A9",X"E5",X"E9",X"A0",X"00",X"00",X"00",X"00",X"9E",X"54",X"5E",
		X"90",X"00",X"00",X"00",X"00",X"9E",X"45",X"5E",X"90",X"00",X"00",X"00",X"00",X"9E",X"5E",X"5E",
		X"90",X"00",X"00",X"00",X"00",X"90",X"E5",X"E0",X"90",X"00",X"00",X"00",X"00",X"80",X"9E",X"90",
		X"80",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"90",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"A9",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"9A",X"90",
		X"00",X"00",X"00",X"00",X"00",X"08",X"90",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"09",X"00",
		X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"A0",X"90",X"00",X"00",X"00",X"00",X"00",X"0A",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E5",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",
		X"00",X"00",X"00",X"09",X"90",X"00",X"94",X"90",X"00",X"00",X"00",X"98",X"00",X"00",X"09",X"00",
		X"00",X"99",X"90",X"00",X"00",X"A9",X"55",X"59",X"A0",X"09",X"80",X"00",X"00",X"9E",X"54",X"5E",
		X"90",X"00",X"00",X"00",X"00",X"0E",X"45",X"4E",X"00",X"00",X"00",X"09",X"00",X"0E",X"44",X"5E",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"54",X"5E",X"90",X"09",X"00",X"00",X"00",X"00",X"95",X"90",
		X"00",X"09",X"90",X"00",X"89",X"90",X"0E",X"90",X"00",X"00",X"80",X"00",X"09",X"00",X"99",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",
		X"80",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"0A",X"A0",X"00",X"07",X"77",X"00",X"00",X"77",X"07",X"00",X"00",X"77",X"77",X"22",X"00",X"07",
		X"74",X"02",X"00",X"03",X"04",X"00",X"00",X"00",X"BB",X"00",X"0B",X"22",X"B0",X"0B",X"22",X"B0",
		X"00",X"BB",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"28",X"43",X"29",X"20",X"31",X"39",
		X"38",X"34",X"2C",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",
		X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"00",X"00",X"00",
		X"A9",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"99",X"00",X"00",X"00",X"00",X"00",X"99",
		X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"0A",X"99",X"98",X"00",X"00",X"00",X"00",X"00",X"09",
		X"98",X"88",X"80",X"00",X"00",X"00",X"00",X"0A",X"98",X"89",X"00",X"00",X"00",X"00",X"00",X"09",
		X"98",X"88",X"00",X"00",X"00",X"00",X"00",X"99",X"9C",X"00",X"00",X"00",X"00",X"00",X"09",X"99",
		X"99",X"C0",X"00",X"00",X"00",X"00",X"99",X"99",X"99",X"E0",X"00",X"00",X"00",X"09",X"99",X"00",
		X"99",X"80",X"00",X"00",X"00",X"09",X"90",X"0A",X"99",X"90",X"00",X"00",X"00",X"09",X"99",X"09",
		X"99",X"90",X"00",X"00",X"00",X"00",X"C8",X"8A",X"99",X"90",X"90",X"00",X"00",X"00",X"08",X"8A",
		X"99",X"90",X"99",X"80",X"00",X"00",X"09",X"09",X"A9",X"90",X"09",X"90",X"00",X"00",X"99",X"99",
		X"80",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"89",X"00",X"00",X"00",X"00",X"00",X"99",X"99",
		X"89",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"90",X"00",X"00",X"00",X"00",X"0A",X"99",
		X"09",X"9A",X"00",X"00",X"00",X"00",X"09",X"90",X"00",X"99",X"00",X"00",X"00",X"0A",X"99",X"00",
		X"00",X"A9",X"90",X"00",X"00",X"99",X"A0",X"00",X"00",X"09",X"90",X"99",X"00",X"09",X"00",X"00",
		X"00",X"00",X"99",X"A0",X"00",X"09",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"A9",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"99",X"00",X"00",X"00",X"00",X"00",X"99",
		X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"0A",X"99",X"98",X"00",X"00",X"00",X"00",X"00",X"09",
		X"98",X"88",X"80",X"00",X"00",X"00",X"00",X"0A",X"98",X"89",X"00",X"00",X"00",X"00",X"00",X"00",
		X"98",X"88",X"00",X"00",X"00",X"00",X"00",X"09",X"8C",X"00",X"00",X"00",X"00",X"00",X"00",X"99",
		X"99",X"C0",X"00",X"00",X"00",X"00",X"09",X"99",X"99",X"E0",X"00",X"00",X"00",X"00",X"99",X"90",
		X"99",X"80",X"00",X"00",X"00",X"00",X"99",X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"99",X"09",
		X"99",X"90",X"00",X"00",X"00",X"00",X"99",X"99",X"99",X"90",X"00",X"00",X"00",X"00",X"CC",X"88",
		X"99",X"90",X"00",X"00",X"00",X"00",X"09",X"88",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"90",
		X"90",X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"98",X"00",X"00",X"00",X"00",X"00",X"09",X"99",
		X"98",X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"98",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A9",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"99",X"00",X"00",X"00",X"00",X"00",X"99",
		X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"0A",X"99",X"98",X"00",X"00",X"00",X"00",X"00",X"09",
		X"98",X"88",X"80",X"00",X"00",X"00",X"00",X"0A",X"98",X"89",X"00",X"00",X"00",X"00",X"00",X"00",
		X"98",X"88",X"00",X"00",X"00",X"00",X"00",X"09",X"8C",X"00",X"00",X"00",X"00",X"00",X"00",X"99",
		X"99",X"C0",X"00",X"00",X"00",X"00",X"09",X"99",X"99",X"E0",X"00",X"00",X"00",X"00",X"99",X"90",
		X"99",X"80",X"00",X"00",X"00",X"00",X"99",X"0A",X"99",X"90",X"00",X"00",X"00",X"00",X"A9",X"99",
		X"99",X"90",X"00",X"00",X"00",X"00",X"09",X"C8",X"8A",X"90",X"00",X"00",X"00",X"00",X"00",X"98",
		X"8A",X"90",X"00",X"00",X"00",X"00",X"00",X"09",X"A9",X"90",X"00",X"00",X"00",X"00",X"00",X"99",
		X"99",X"80",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"80",X"00",X"00",X"00",X"00",X"00",X"99",
		X"99",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"99",
		X"AA",X"00",X"00",X"00",X"00",X"00",X"09",X"90",X"A9",X"A0",X"00",X"00",X"00",X"0A",X"99",X"00",
		X"0A",X"90",X"00",X"00",X"00",X"99",X"90",X"00",X"0A",X"90",X"00",X"00",X"00",X"09",X"00",X"00",
		X"0A",X"A0",X"00",X"00",X"00",X"09",X"90",X"00",X"09",X"09",X"90",X"00",X"00",X"00",X"00",X"09",
		X"9A",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"AA",X"00",X"00",X"00",X"00",X"00",X"99",X"99",
		X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"89",X"99",X"A0",X"00",X"00",X"00",X"00",X"08",X"88",
		X"89",X"90",X"00",X"00",X"00",X"00",X"00",X"98",X"89",X"A0",X"00",X"00",X"00",X"00",X"00",X"88",
		X"89",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"C9",X"99",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"99",X"99",X"90",X"00",X"00",X"00",X"00",X"0E",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"08",
		X"99",X"00",X"99",X"90",X"00",X"00",X"00",X"09",X"99",X"A0",X"09",X"90",X"00",X"00",X"00",X"09",
		X"99",X"90",X"99",X"90",X"00",X"00",X"09",X"09",X"99",X"A8",X"8C",X"00",X"00",X"08",X"99",X"09",
		X"99",X"A8",X"80",X"00",X"00",X"09",X"90",X"09",X"9A",X"90",X"90",X"00",X"00",X"00",X"00",X"00",
		X"08",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"98",X"99",X"99",X"00",X"00",X"00",X"00",X"0A",
		X"98",X"99",X"99",X"00",X"00",X"00",X"00",X"09",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"A9",
		X"90",X"99",X"A0",X"00",X"00",X"00",X"00",X"99",X"00",X"09",X"90",X"00",X"00",X"00",X"09",X"9A",
		X"00",X"00",X"99",X"A0",X"00",X"99",X"09",X"90",X"00",X"00",X"0A",X"99",X"00",X"0A",X"99",X"00",
		X"00",X"00",X"00",X"90",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"00",X"09",
		X"9A",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"AA",X"00",X"00",X"00",X"00",X"00",X"99",X"99",
		X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"89",X"99",X"A0",X"00",X"00",X"00",X"00",X"08",X"88",
		X"89",X"90",X"00",X"00",X"00",X"00",X"00",X"98",X"89",X"A0",X"00",X"00",X"00",X"00",X"00",X"88",
		X"89",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C8",X"90",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"0E",X"99",X"99",X"90",X"00",X"00",X"00",X"00",X"08",
		X"99",X"09",X"99",X"00",X"00",X"00",X"00",X"09",X"99",X"00",X"99",X"00",X"00",X"00",X"00",X"09",
		X"99",X"90",X"99",X"00",X"00",X"00",X"00",X"09",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"09",
		X"99",X"88",X"CC",X"00",X"00",X"00",X"00",X"09",X"99",X"88",X"90",X"00",X"00",X"00",X"00",X"00",
		X"09",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"89",X"99",X"90",X"00",X"00",X"00",X"00",X"00",
		X"89",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"89",X"99",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"AA",X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"09",X"00",X"00",X"00",X"00",X"00",X"09",
		X"9A",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"AA",X"00",X"00",X"00",X"00",X"00",X"99",X"99",
		X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"89",X"99",X"A0",X"00",X"00",X"00",X"00",X"08",X"88",
		X"89",X"90",X"00",X"00",X"00",X"00",X"00",X"98",X"89",X"A0",X"00",X"00",X"00",X"00",X"00",X"88",
		X"89",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C8",X"90",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"0E",X"99",X"99",X"90",X"00",X"00",X"00",X"00",X"08",
		X"99",X"09",X"99",X"00",X"00",X"00",X"00",X"09",X"99",X"A0",X"99",X"00",X"00",X"00",X"00",X"09",
		X"99",X"99",X"9A",X"00",X"00",X"00",X"00",X"09",X"A8",X"8C",X"90",X"00",X"00",X"00",X"00",X"09",
		X"A8",X"89",X"00",X"00",X"00",X"00",X"00",X"09",X"9A",X"90",X"00",X"00",X"00",X"00",X"00",X"08",
		X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"08",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"08",
		X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"99",X"A0",X"00",X"00",X"00",X"00",X"0A",X"9A",X"09",X"90",X"00",X"00",X"00",X"00",X"09",
		X"A0",X"00",X"99",X"A0",X"00",X"00",X"00",X"09",X"A0",X"00",X"09",X"99",X"00",X"00",X"00",X"0A",
		X"A0",X"00",X"00",X"90",X"00",X"00",X"09",X"90",X"90",X"00",X"09",X"90",X"00",X"00",X"00",X"0A",
		X"9A",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"00",X"00",X"09",X"99",
		X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"89",
		X"89",X"80",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"08",
		X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"89",X"00",X"00",X"00",X"00",X"00",X"A9",X"9C",
		X"5C",X"99",X"A0",X"00",X"00",X"00",X"99",X"98",X"58",X"99",X"90",X"00",X"00",X"00",X"9A",X"99",
		X"C9",X"9A",X"90",X"00",X"00",X"00",X"9A",X"99",X"89",X"9A",X"90",X"00",X"00",X"00",X"9A",X"99",
		X"A9",X"9A",X"90",X"00",X"00",X"00",X"AA",X"99",X"A9",X"9A",X"A0",X"00",X"00",X"00",X"90",X"99",
		X"A9",X"99",X"90",X"00",X"00",X"00",X"80",X"99",X"A9",X"98",X"80",X"00",X"00",X"00",X"00",X"AA",
		X"AA",X"A9",X"80",X"00",X"00",X"00",X"00",X"09",X"A9",X"09",X"90",X"00",X"00",X"00",X"00",X"09",
		X"A9",X"09",X"90",X"00",X"00",X"00",X"00",X"09",X"A9",X"09",X"90",X"00",X"00",X"00",X"00",X"09",
		X"A9",X"09",X"90",X"00",X"00",X"00",X"00",X"09",X"A9",X"00",X"00",X"00",X"00",X"00",X"00",X"09",
		X"A9",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"A9",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",
		X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"99",X"A9",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"99",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"98",X"98",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"99",
		X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"98",X"90",X"00",X"00",X"00",X"00",X"00",X"0A",X"99",X"E5",X"E9",X"9A",X"00",X"00",X"00",
		X"00",X"09",X"9E",X"55",X"5E",X"99",X"00",X"00",X"00",X"00",X"09",X"A5",X"55",X"55",X"A9",X"00",
		X"00",X"00",X"00",X"09",X"A5",X"55",X"55",X"A9",X"00",X"00",X"00",X"00",X"09",X"A5",X"55",X"55",
		X"A9",X"00",X"00",X"00",X"00",X"0A",X"AE",X"5E",X"5E",X"AA",X"00",X"00",X"00",X"00",X"09",X"A9",
		X"EE",X"E9",X"99",X"00",X"00",X"00",X"00",X"08",X"09",X"9A",X"99",X"88",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"AA",X"AA",X"98",X"00",X"00",X"00",X"00",X"00",X"00",X"9A",X"90",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"9A",X"90",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"9A",X"90",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"9A",X"90",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"9A",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9A",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"9A",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"AA",X"AA",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"9A",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A9",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"99",
		X"90",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"09",X"E5",X"E9",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"90",X"98",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"95",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"84",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"99",X"E5",X"E9",X"9A",X"00",X"00",X"00",X"00",X"09",X"EE",X"55",
		X"4E",X"E9",X"00",X"00",X"00",X"00",X"09",X"A5",X"55",X"55",X"A9",X"00",X"00",X"00",X"00",X"09",
		X"A4",X"55",X"54",X"A9",X"00",X"00",X"00",X"00",X"09",X"A5",X"45",X"55",X"A9",X"00",X"00",X"00",
		X"00",X"0A",X"AE",X"5E",X"5E",X"AA",X"00",X"00",X"00",X"00",X"09",X"09",X"E4",X"E9",X"99",X"00",
		X"00",X"00",X"00",X"08",X"09",X"95",X"99",X"88",X"00",X"00",X"00",X"00",X"00",X"0A",X"A0",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"A0",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"90",
		X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"98",X"00",X"00",X"00",
		X"00",X"00",X"90",X"90",X"90",X"99",X"90",X"00",X"00",X"00",X"09",X"00",X"90",X"99",X"00",X"00",
		X"00",X"00",X"00",X"99",X"09",X"E5",X"E9",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"95",X"99",X"00",X"00",X"00",X"00",X"09",X"90",X"00",
		X"84",X"80",X"09",X"98",X"00",X"00",X"09",X"80",X"00",X"90",X"90",X"00",X"88",X"00",X"00",X"00",
		X"00",X"00",X"E5",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"55",X"4E",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"A5",X"55",X"55",X"A0",X"00",X"00",X"00",X"80",X"00",X"A4",X"54",X"54",X"A0",
		X"99",X"00",X"00",X"00",X"00",X"05",X"45",X"55",X"A0",X"09",X"90",X"00",X"00",X"00",X"0E",X"5E",
		X"5E",X"00",X"00",X"90",X"00",X"00",X"88",X"09",X"E4",X"E9",X"00",X"00",X"00",X"00",X"09",X"90",
		X"09",X"05",X"99",X"00",X"00",X"00",X"00",X"09",X"90",X"0A",X"00",X"AA",X"00",X"90",X"00",X"00",
		X"00",X"00",X"09",X"00",X"90",X"09",X"90",X"00",X"00",X"00",X"00",X"09",X"00",X"90",X"00",X"08",
		X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"90",
		X"00",X"09",X"09",X"80",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"09",X"90",X"00",X"00",X"00",X"09",X"90",X"00",X"00",X"09",X"90",X"00",X"00",X"00",X"09",X"90",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"09",X"9A",X"00",X"00",X"00",X"00",X"09",
		X"99",X"99",X"9A",X"00",X"00",X"00",X"00",X"08",X"99",X"A0",X"00",X"00",X"00",X"00",X"88",X"89",
		X"A0",X"00",X"00",X"00",X"00",X"08",X"89",X"A0",X"00",X"00",X"00",X"00",X"00",X"0C",X"99",X"00",
		X"00",X"00",X"00",X"00",X"C9",X"99",X"90",X"00",X"00",X"00",X"00",X"E9",X"9A",X"99",X"00",X"00",
		X"00",X"00",X"89",X"A0",X"A9",X"90",X"00",X"00",X"0A",X"99",X"90",X"A9",X"90",X"00",X"00",X"9A",
		X"99",X"9A",X"99",X"00",X"00",X"08",X"90",X"99",X"A8",X"8C",X"00",X"00",X"09",X"00",X"99",X"AA",
		X"90",X"00",X"00",X"00",X"00",X"00",X"89",X"99",X"00",X"00",X"00",X"00",X"A9",X"89",X"99",X"00",
		X"00",X"00",X"00",X"99",X"89",X"99",X"00",X"00",X"00",X"0A",X"9A",X"0A",X"00",X"00",X"00",X"00",
		X"A9",X"A0",X"09",X"90",X"00",X"00",X"90",X"99",X"00",X"00",X"99",X"A0",X"00",X"A9",X"9A",X"00",
		X"00",X"00",X"99",X"00",X"0A",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"00",X"00",X"09",X"9A",X"00",X"00",X"00",X"00",X"09",X"99",X"99",X"9A",X"00",X"00",X"00",
		X"00",X"08",X"99",X"A0",X"00",X"00",X"00",X"00",X"88",X"89",X"A0",X"00",X"00",X"00",X"00",X"08",
		X"89",X"A0",X"00",X"00",X"00",X"00",X"00",X"0C",X"90",X"00",X"00",X"00",X"00",X"00",X"C9",X"9A",
		X"00",X"00",X"00",X"00",X"00",X"E9",X"99",X"A0",X"00",X"00",X"00",X"00",X"89",X"A9",X"9A",X"00",
		X"00",X"00",X"00",X"99",X"A0",X"99",X"00",X"00",X"00",X"00",X"99",X"90",X"99",X"00",X"00",X"00",
		X"00",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"99",X"88",X"C0",X"00",X"00",X"00",X"00",X"0A",
		X"A9",X"00",X"00",X"00",X"00",X"00",X"08",X"99",X"90",X"00",X"00",X"00",X"00",X"08",X"99",X"90",
		X"00",X"00",X"00",X"00",X"08",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"99",X"A9",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"09",X"9A",X"00",
		X"00",X"00",X"00",X"09",X"99",X"99",X"9A",X"00",X"00",X"00",X"00",X"08",X"99",X"A0",X"00",X"00",
		X"00",X"00",X"88",X"89",X"A0",X"00",X"00",X"00",X"00",X"08",X"89",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"90",X"00",X"00",X"00",X"00",X"00",X"C9",X"99",X"00",X"00",X"00",X"00",X"00",X"E9",
		X"99",X"90",X"00",X"00",X"00",X"00",X"89",X"0A",X"99",X"00",X"00",X"00",X"0A",X"99",X"90",X"99",
		X"00",X"00",X"00",X"00",X"99",X"99",X"90",X"00",X"00",X"00",X"00",X"98",X"8C",X"00",X"00",X"00",
		X"00",X"00",X"9A",X"90",X"00",X"00",X"00",X"00",X"00",X"89",X"99",X"00",X"00",X"00",X"00",X"00",
		X"89",X"99",X"00",X"00",X"00",X"00",X"00",X"89",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"A9",X"90",X"00",X"00",X"00",X"00",X"9A",X"00",X"99",X"A0",
		X"00",X"00",X"00",X"9A",X"00",X"00",X"99",X"00",X"00",X"99",X"A9",X"00",X"09",X"90",X"00",X"00",
		X"00",X"0A",X"A0",X"00",X"00",X"00",X"00",X"00",X"09",X"9A",X"00",X"00",X"00",X"00",X"00",X"99",
		X"99",X"90",X"00",X"00",X"00",X"00",X"0A",X"AA",X"00",X"00",X"00",X"00",X"00",X"09",X"89",X"00",
		X"00",X"00",X"00",X"00",X"08",X"98",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",
		X"00",X"0A",X"9C",X"58",X"9A",X"00",X"00",X"00",X"09",X"99",X"E9",X"99",X"00",X"00",X"00",X"09",
		X"09",X"89",X"09",X"00",X"00",X"00",X"09",X"A9",X"99",X"A9",X"00",X"00",X"00",X"09",X"99",X"A9",
		X"99",X"00",X"00",X"00",X"0A",X"99",X"A9",X"9A",X"00",X"00",X"00",X"08",X"99",X"A9",X"98",X"00",
		X"00",X"00",X"00",X"0A",X"AA",X"0A",X"A0",X"00",X"00",X"00",X"09",X"A9",X"09",X"A0",X"00",X"00",
		X"00",X"09",X"A9",X"09",X"A0",X"00",X"00",X"00",X"09",X"A9",X"09",X"A0",X"00",X"00",X"00",X"09",
		X"A9",X"00",X"00",X"00",X"00",X"00",X"09",X"A9",X"00",X"00",X"00",X"00",X"00",X"A9",X"99",X"A0",
		X"00",X"00",X"00",X"00",X"99",X"09",X"90",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"A9",X"90",X"00",X"00",X"00",X"00",X"A9",X"99",X"99",X"90",X"00",X"00",X"00",
		X"0A",X"99",X"80",X"00",X"00",X"00",X"00",X"0A",X"98",X"88",X"00",X"00",X"00",X"00",X"0A",X"98",
		X"80",X"00",X"00",X"00",X"00",X"99",X"C0",X"00",X"00",X"00",X"00",X"09",X"99",X"9C",X"00",X"00",
		X"00",X"00",X"99",X"A9",X"9E",X"00",X"00",X"00",X"09",X"9A",X"0A",X"98",X"00",X"00",X"00",X"09",
		X"9A",X"09",X"99",X"A0",X"00",X"00",X"00",X"99",X"A9",X"99",X"A9",X"00",X"00",X"00",X"C8",X"8A",
		X"99",X"09",X"80",X"00",X"00",X"09",X"AA",X"99",X"00",X"90",X"00",X"00",X"99",X"98",X"00",X"00",
		X"00",X"00",X"00",X"99",X"98",X"9A",X"00",X"00",X"00",X"00",X"99",X"98",X"99",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"A9",X"A0",X"00",X"00",X"00",X"09",X"90",X"0A",X"9A",X"00",X"00",X"0A",X"99",
		X"00",X"00",X"99",X"09",X"00",X"99",X"00",X"00",X"00",X"A9",X"9A",X"00",X"09",X"99",X"00",X"00",
		X"09",X"A0",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"A9",X"90",X"00",
		X"00",X"00",X"00",X"A9",X"99",X"99",X"90",X"00",X"00",X"00",X"0A",X"99",X"80",X"00",X"00",X"00",
		X"00",X"0A",X"98",X"88",X"00",X"00",X"00",X"00",X"0A",X"98",X"80",X"00",X"00",X"00",X"00",X"09",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"A9",X"9C",X"00",X"00",X"00",X"00",X"0A",X"99",X"9E",X"00",
		X"00",X"00",X"00",X"A9",X"9A",X"98",X"00",X"00",X"00",X"00",X"99",X"0A",X"99",X"00",X"00",X"00",
		X"00",X"99",X"09",X"99",X"00",X"00",X"00",X"00",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"0C",
		X"88",X"99",X"00",X"00",X"00",X"00",X"00",X"9A",X"A0",X"00",X"00",X"00",X"00",X"09",X"99",X"80",
		X"00",X"00",X"00",X"00",X"09",X"99",X"80",X"00",X"00",X"00",X"00",X"09",X"99",X"80",X"00",X"00",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"9A",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"A9",X"90",X"00",X"00",X"00",X"00",X"A9",X"99",X"99",
		X"90",X"00",X"00",X"00",X"0A",X"99",X"80",X"00",X"00",X"00",X"00",X"0A",X"98",X"88",X"00",X"00",
		X"00",X"00",X"0A",X"98",X"80",X"00",X"00",X"00",X"00",X"09",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"99",X"9C",X"00",X"00",X"00",X"00",X"09",X"99",X"9E",X"00",X"00",X"00",X"00",X"99",X"A0",X"98",
		X"00",X"00",X"00",X"00",X"99",X"09",X"99",X"A0",X"00",X"00",X"00",X"09",X"99",X"99",X"00",X"00",
		X"00",X"00",X"00",X"C8",X"89",X"00",X"00",X"00",X"00",X"00",X"09",X"A9",X"00",X"00",X"00",X"00",
		X"00",X"99",X"98",X"00",X"00",X"00",X"00",X"00",X"99",X"98",X"00",X"00",X"00",X"00",X"00",X"99",
		X"98",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"09",X"9A",X"A0",X"00",
		X"00",X"00",X"0A",X"99",X"00",X"A9",X"00",X"00",X"00",X"99",X"00",X"00",X"A9",X"00",X"00",X"00",
		X"09",X"90",X"00",X"9A",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"98",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"89",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"A9",X"95",X"99",X"A0",X"00",X"00",X"00",X"00",X"00",X"99",X"E5",X"E9",X"90",
		X"00",X"00",X"00",X"00",X"00",X"9E",X"55",X"5E",X"90",X"00",X"00",X"00",X"00",X"00",X"9E",X"55",
		X"5E",X"90",X"00",X"00",X"00",X"00",X"00",X"9E",X"55",X"5E",X"90",X"00",X"00",X"00",X"00",X"00",
		X"A9",X"E5",X"E9",X"A0",X"00",X"00",X"00",X"00",X"00",X"89",X"9A",X"99",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"AA",X"A0",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"9A",X"90",X"9A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"9A",X"90",X"9A",X"00",X"00",X"00",X"00",X"00",X"00",X"9A",X"90",
		X"9A",X"00",X"00",X"00",X"00",X"00",X"00",X"9A",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"9A",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"99",X"9A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"90",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",
		X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"E5",X"E9",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"A0",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"95",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"84",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"A9",X"E5",X"E9",X"A0",X"00",X"00",X"00",X"00",X"00",X"9E",X"54",X"5E",
		X"90",X"00",X"00",X"00",X"00",X"00",X"95",X"55",X"45",X"90",X"00",X"00",X"00",X"00",X"00",X"95",
		X"45",X"55",X"90",X"00",X"00",X"00",X"00",X"00",X"9E",X"45",X"5E",X"90",X"00",X"00",X"00",X"00",
		X"00",X"AE",X"E5",X"EE",X"A0",X"00",X"00",X"00",X"00",X"00",X"89",X"E5",X"E9",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9A",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"9A",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9A",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9A",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"9A",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"99",X"9A",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"90",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"98",X"00",X"00",X"00",X"00",X"09",X"00",X"A0",X"A0",X"99",X"00",X"00",X"00",X"00",X"09",X"90",
		X"90",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"E5",X"E9",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"A0",X"AE",X"00",X"00",X"00",X"00",X"09",X"90",X"00",X"95",X"90",X"00",X"99",X"90",
		X"00",X"09",X"80",X"00",X"84",X"80",X"00",X"09",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"5E",X"E5",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",X"9E",X"54",
		X"5E",X"90",X"00",X"00",X"00",X"00",X"00",X"95",X"55",X"45",X"A0",X"00",X"00",X"00",X"80",X"00",
		X"A5",X"45",X"55",X"A0",X"09",X"00",X"00",X"00",X"00",X"0E",X"44",X"55",X"A0",X"00",X"99",X"00",
		X"00",X"00",X"0E",X"E4",X"EE",X"00",X"00",X"09",X"00",X"00",X"80",X"09",X"E5",X"E9",X"00",X"00",
		X"00",X"00",X"09",X"90",X"00",X"AE",X"A0",X"00",X"90",X"00",X"00",X"09",X"90",X"00",X"90",X"09",
		X"09",X"90",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"09",X"80",X"00",X"00",X"90",X"98",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"09",X"90",X"00",X"00",X"0F",X"88",X"F0",X"00",X"00",
		X"00",X"00",X"F8",X"86",X"9F",X"00",X"00",X"00",X"00",X"F8",X"66",X"9F",X"00",X"00",X"00",X"00",
		X"F9",X"99",X"AF",X"00",X"00",X"00",X"0F",X"88",X"88",X"89",X"F0",X"00",X"00",X"0F",X"9A",X"AA",
		X"A9",X"FF",X"00",X"00",X"00",X"FB",X"97",X"7C",X"77",X"00",X"00",X"0F",X"75",X"B5",X"7F",X"78",
		X"F0",X"00",X"0F",X"5F",X"95",X"5F",X"88",X"8F",X"00",X"0F",X"F9",X"88",X"88",X"88",X"F0",X"00",
		X"F8",X"98",X"88",X"69",X"8F",X"00",X"00",X"89",X"A8",X"86",X"FC",X"8F",X"00",X"00",X"87",X"79",
		X"88",X"C8",X"AF",X"00",X"00",X"FB",X"B9",X"88",X"88",X"AF",X"00",X"00",X"0F",X"88",X"88",X"88",
		X"AF",X"00",X"00",X"00",X"F9",X"99",X"9F",X"F0",X"00",X"00",X"FC",X"FF",X"A8",X"F0",X"00",X"00",
		X"00",X"FE",X"99",X"98",X"F0",X"00",X"00",X"00",X"0F",X"EE",X"E8",X"F0",X"00",X"00",X"00",X"00",
		X"FF",X"F8",X"FF",X"F0",X"00",X"00",X"00",X"00",X"F8",X"88",X"CF",X"00",X"00",X"00",X"00",X"FE",
		X"EE",X"EF",X"00",X"00",X"00",X"0F",X"88",X"F0",X"00",X"00",X"00",X"00",X"F8",X"86",X"9F",X"00",
		X"00",X"00",X"00",X"F8",X"66",X"95",X"F0",X"00",X"00",X"00",X"F9",X"99",X"9C",X"5F",X"00",X"00",
		X"0F",X"88",X"88",X"89",X"C5",X"F0",X"00",X"0F",X"9A",X"AA",X"A9",X"FC",X"7F",X"00",X"00",X"FB",
		X"F7",X"7F",X"F7",X"2F",X"00",X"0F",X"75",X"B5",X"7F",X"F8",X"8F",X"00",X"0F",X"5F",X"A5",X"5F",
		X"F8",X"8F",X"00",X"00",X"F9",X"88",X"88",X"88",X"8F",X"00",X"0F",X"88",X"88",X"68",X"88",X"F0",
		X"00",X"08",X"98",X"86",X"FC",X"8F",X"00",X"00",X"08",X"99",X"88",X"C8",X"9F",X"00",X"00",X"08",
		X"77",X"88",X"88",X"9F",X"00",X"00",X"0F",X"BB",X"88",X"88",X"9F",X"00",X"00",X"00",X"F9",X"99",
		X"9F",X"F0",X"00",X"00",X"00",X"0F",X"98",X"F0",X"00",X"00",X"00",X"00",X"0F",X"98",X"F0",X"00",
		X"00",X"00",X"0F",X"0F",X"98",X"F0",X"00",X"00",X"00",X"FC",X"FF",X"98",X"FF",X"F0",X"00",X"00",
		X"FE",X"99",X"98",X"88",X"CF",X"00",X"00",X"0F",X"EE",X"EE",X"EE",X"F0",X"00",X"00",X"00",X"0F",
		X"88",X"F0",X"00",X"C4",X"00",X"00",X"F8",X"86",X"9F",X"0F",X"C5",X"F0",X"00",X"F8",X"66",X"9F",
		X"0F",X"C5",X"F0",X"00",X"F9",X"99",X"AF",X"0F",X"C5",X"F0",X"0F",X"88",X"88",X"89",X"FF",X"C5",
		X"F0",X"0F",X"9A",X"AA",X"A9",X"FF",X"77",X"F0",X"00",X"FB",X"97",X"7F",X"08",X"72",X"F0",X"0F",
		X"75",X"B5",X"7F",X"F8",X"87",X"F0",X"0F",X"5F",X"95",X"5F",X"88",X"8F",X"00",X"0F",X"F9",X"88",
		X"88",X"88",X"F0",X"00",X"F9",X"88",X"88",X"69",X"8F",X"00",X"00",X"87",X"79",X"86",X"FC",X"8F",
		X"00",X"00",X"8B",X"B9",X"88",X"C8",X"AF",X"00",X"00",X"F9",X"98",X"88",X"88",X"AF",X"00",X"00",
		X"0F",X"88",X"88",X"88",X"AF",X"00",X"00",X"00",X"F9",X"99",X"9F",X"F0",X"00",X"00",X"00",X"FF",
		X"A8",X"FF",X"CF",X"00",X"00",X"00",X"0F",X"98",X"88",X"EF",X"00",X"00",X"00",X"0F",X"9E",X"EE",
		X"F0",X"00",X"00",X"0F",X"FF",X"9F",X"00",X"00",X"00",X"00",X"FC",X"99",X"9F",X"00",X"00",X"00",
		X"00",X"0E",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"8F",X"00",X"00",X"00",
		X"00",X"0F",X"96",X"88",X"F0",X"00",X"00",X"00",X"0F",X"96",X"68",X"F0",X"00",X"00",X"00",X"0F",
		X"A9",X"99",X"F0",X"00",X"00",X"00",X"F9",X"88",X"88",X"8F",X"00",X"00",X"0F",X"F9",X"AA",X"AA",
		X"9F",X"00",X"00",X"07",X"7C",X"77",X"9B",X"F0",X"00",X"00",X"F8",X"7F",X"75",X"B5",X"7F",X"00",
		X"0F",X"88",X"8F",X"55",X"9F",X"5F",X"00",X"00",X"F8",X"88",X"88",X"89",X"FF",X"00",X"00",X"0F",
		X"89",X"68",X"88",X"98",X"F0",X"00",X"0F",X"8C",X"F6",X"88",X"A9",X"80",X"00",X"0F",X"A8",X"C8",
		X"89",X"77",X"80",X"00",X"0F",X"A8",X"88",X"89",X"BB",X"F0",X"00",X"0F",X"A8",X"88",X"88",X"8F",
		X"00",X"00",X"00",X"FF",X"99",X"99",X"F0",X"00",X"00",X"00",X"00",X"F8",X"AF",X"FC",X"F0",X"00",
		X"00",X"00",X"F8",X"99",X"9E",X"F0",X"00",X"00",X"00",X"F8",X"EE",X"EF",X"00",X"00",X"00",X"FF",
		X"F8",X"FF",X"F0",X"00",X"00",X"0F",X"C8",X"88",X"F0",X"00",X"00",X"00",X"0F",X"EE",X"EE",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"F8",X"8F",X"00",X"00",X"00",X"00",X"0F",X"96",X"88",X"F0",X"00",
		X"00",X"00",X"F5",X"96",X"68",X"F0",X"00",X"00",X"0F",X"5C",X"99",X"99",X"F0",X"00",X"00",X"F5",
		X"C9",X"88",X"88",X"8F",X"00",X"0F",X"7C",X"F9",X"AA",X"AA",X"9F",X"00",X"0F",X"27",X"FF",X"77",
		X"FB",X"F0",X"00",X"0F",X"88",X"FF",X"75",X"B5",X"7F",X"00",X"0F",X"88",X"FF",X"55",X"AF",X"5F",
		X"00",X"0F",X"88",X"88",X"88",X"89",X"F0",X"00",X"00",X"F8",X"88",X"68",X"88",X"8F",X"00",X"00",
		X"0F",X"8C",X"F6",X"88",X"98",X"00",X"00",X"0F",X"98",X"C8",X"89",X"98",X"00",X"00",X"0F",X"98",
		X"88",X"87",X"78",X"00",X"00",X"0F",X"98",X"88",X"8B",X"BF",X"00",X"00",X"00",X"FF",X"99",X"99",
		X"F0",X"00",X"00",X"00",X"00",X"F8",X"9F",X"00",X"00",X"00",X"00",X"00",X"F8",X"9F",X"00",X"00",
		X"00",X"00",X"00",X"F8",X"9F",X"0F",X"00",X"00",X"00",X"FF",X"F8",X"9F",X"FC",X"F0",X"00",X"0F",
		X"C8",X"88",X"99",X"9E",X"F0",X"00",X"00",X"FE",X"EE",X"EE",X"EF",X"00",X"04",X"C0",X"00",X"F8",
		X"8F",X"00",X"00",X"F5",X"CF",X"0F",X"96",X"88",X"F0",X"00",X"F5",X"CF",X"0F",X"96",X"68",X"F0",
		X"00",X"F5",X"CF",X"0F",X"A9",X"99",X"F0",X"00",X"F5",X"CF",X"F9",X"88",X"88",X"8F",X"00",X"F7",
		X"7F",X"F9",X"AA",X"AA",X"9F",X"00",X"F2",X"78",X"0F",X"77",X"9B",X"F0",X"00",X"F7",X"88",X"FF",
		X"75",X"B5",X"7F",X"00",X"0F",X"88",X"8F",X"55",X"9F",X"5F",X"00",X"00",X"F8",X"88",X"88",X"89",
		X"FF",X"00",X"00",X"0F",X"89",X"68",X"88",X"89",X"F0",X"00",X"0F",X"8C",X"F6",X"89",X"77",X"80",
		X"00",X"0F",X"A8",X"C8",X"89",X"BB",X"80",X"00",X"0F",X"A8",X"88",X"88",X"99",X"F0",X"00",X"0F",
		X"A8",X"88",X"88",X"8F",X"00",X"00",X"00",X"FF",X"99",X"99",X"F0",X"00",X"00",X"0F",X"CF",X"F8",
		X"AF",X"F0",X"00",X"00",X"0F",X"E8",X"88",X"9F",X"00",X"00",X"00",X"00",X"FE",X"EE",X"9F",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"9F",X"FF",X"00",X"00",X"00",X"00",X"0F",X"99",X"9C",X"F0",X"00",
		X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"50",X"00",X"00",X"00",X"00",
		X"00",X"A6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"88",
		X"E4",X"56",X"D6",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"D6",
		X"C0",X"09",X"8D",X"DD",X"D8",X"64",X"48",X"6D",X"D6",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"66",X"00",X"8D",X"DD",X"DD",X"DD",X"88",X"58",X"86",X"DD",X"DC",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"88",X"D6",X"99",X"98",X"88",X"C6",
		X"88",X"88",X"6D",X"DD",X"6C",X"66",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"DD",X"6D",
		X"99",X"88",X"88",X"99",X"9D",X"D9",X"99",X"98",X"66",X"6C",X"D6",X"50",X"00",X"00",X"00",X"00",
		X"C6",X"DD",X"DD",X"DD",X"D8",X"88",X"89",X"99",X"9F",X"F6",X"68",X"89",X"86",X"66",X"6D",X"DD",
		X"DC",X"00",X"00",X"0C",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"68",X"99",X"FF",X"F9",X"9C",X"CA",
		X"98",X"66",X"DD",X"DD",X"DD",X"DD",X"D4",X"00",X"6D",X"DD",X"DD",X"DD",X"66",X"66",X"6D",X"D6",
		X"68",X"88",X"88",X"CC",X"69",X"86",X"6D",X"DD",X"DD",X"D6",X"66",X"65",X"00",X"DD",X"DD",X"DD",
		X"66",X"DD",X"DD",X"66",X"6D",X"88",X"88",X"88",X"86",X"66",X"6D",X"DD",X"D6",X"66",X"66",X"6C",
		X"00",X"00",X"C6",X"DD",X"D6",X"6D",X"DD",X"DD",X"DD",X"6C",X"88",X"82",X"28",X"88",X"DD",X"DD",
		X"66",X"66",X"66",X"6C",X"00",X"00",X"00",X"00",X"44",X"44",X"DD",X"D6",X"66",X"6D",X"D6",X"C9",
		X"99",X"99",X"99",X"66",X"66",X"66",X"6C",X"CC",X"6C",X"6C",X"00",X"00",X"00",X"05",X"4C",X"DD",
		X"66",X"66",X"66",X"DD",X"6C",X"99",X"99",X"99",X"96",X"6C",X"90",X"00",X"09",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"8D",X"66",X"66",X"66",X"66",X"D6",X"00",X"00",X"00",X"00",X"09",X"98",
		X"DC",X"89",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"98",X"89",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"98",X"88",X"99",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A9",
		X"9A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A9",X"99",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",
		X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"4E",X"00",X"00",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"88",X"5E",X"56",X"D6",X"00",X"00",X"00",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"C0",X"09",X"8D",X"DD",X"D8",X"65",
		X"58",X"6D",X"D6",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C6",X"00",
		X"8D",X"DD",X"DD",X"DD",X"88",X"E8",X"86",X"DD",X"DC",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"88",X"D6",X"99",X"98",X"88",X"C6",X"88",X"88",X"6D",X"DD",X"6C",X"66",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"DD",X"6D",X"99",X"88",X"88",X"99",X"9D",X"D9",
		X"99",X"98",X"66",X"6C",X"D6",X"50",X"00",X"00",X"00",X"00",X"C6",X"DD",X"DD",X"DD",X"D8",X"88",
		X"89",X"99",X"9F",X"F6",X"68",X"89",X"86",X"66",X"6D",X"DD",X"DC",X"00",X"00",X"0C",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"68",X"99",X"FF",X"F9",X"9C",X"CA",X"98",X"66",X"DD",X"DD",X"DD",X"DD",
		X"D4",X"00",X"6D",X"DD",X"DD",X"DD",X"66",X"66",X"6D",X"D6",X"68",X"88",X"88",X"CC",X"69",X"86",
		X"6D",X"DD",X"DD",X"D6",X"66",X"65",X"00",X"DD",X"DD",X"DD",X"66",X"DD",X"DD",X"66",X"6D",X"88",
		X"88",X"88",X"86",X"66",X"6D",X"DD",X"D6",X"66",X"66",X"6C",X"00",X"00",X"C6",X"DD",X"D6",X"6D",
		X"DD",X"DD",X"DD",X"6C",X"88",X"82",X"28",X"88",X"DD",X"DD",X"66",X"66",X"66",X"6C",X"00",X"00",
		X"00",X"00",X"E5",X"55",X"DD",X"D6",X"66",X"6D",X"D6",X"C9",X"99",X"99",X"99",X"66",X"66",X"66",
		X"6C",X"CC",X"66",X"C0",X"00",X"00",X"00",X"0E",X"5C",X"DD",X"66",X"66",X"66",X"DD",X"6C",X"99",
		X"99",X"99",X"96",X"6C",X"90",X"00",X"09",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"8D",X"66",
		X"66",X"66",X"66",X"D6",X"00",X"00",X"00",X"00",X"09",X"98",X"DC",X"89",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"98",X"89",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"98",X"88",
		X"99",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A9",X"9A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"A9",X"99",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"6A",X"00",X"00",X"00",X"00",X"00",X"05",X"50",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"6D",
		X"65",X"4E",X"88",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"00",X"6D",X"D6",X"84",X"46",X"8D",X"DD",X"D8",X"90",X"0C",X"6D",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"CD",X"DD",X"68",X"85",X"88",X"DD",X"DD",X"DD",X"D8",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"66",X"C6",X"DD",X"D6",X"88",X"88",
		X"6C",X"88",X"89",X"99",X"6D",X"88",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"6D",
		X"C6",X"66",X"89",X"99",X"9D",X"D9",X"99",X"88",X"88",X"99",X"D6",X"DD",X"66",X"00",X"00",X"00",
		X"00",X"00",X"00",X"CD",X"DD",X"D6",X"66",X"68",X"98",X"86",X"6F",X"F9",X"99",X"98",X"88",X"8D",
		X"DD",X"DD",X"DD",X"6C",X"00",X"00",X"00",X"4D",X"DD",X"DD",X"DD",X"DD",X"66",X"89",X"AC",X"C9",
		X"9F",X"FF",X"99",X"86",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"C0",X"00",X"56",X"66",X"6D",X"DD",
		X"DD",X"D6",X"68",X"96",X"CC",X"88",X"88",X"86",X"6D",X"D6",X"66",X"66",X"DD",X"DD",X"DD",X"D6",
		X"00",X"00",X"C6",X"66",X"66",X"6D",X"DD",X"D6",X"66",X"68",X"88",X"88",X"88",X"D6",X"66",X"DD",
		X"DD",X"66",X"DD",X"DD",X"DD",X"00",X"00",X"00",X"C6",X"66",X"66",X"66",X"DD",X"DD",X"88",X"82",
		X"28",X"88",X"C6",X"DD",X"DD",X"DD",X"D6",X"6D",X"DD",X"6C",X"00",X"00",X"C6",X"C6",X"CC",X"C6",
		X"66",X"66",X"66",X"99",X"99",X"99",X"9C",X"6D",X"D6",X"66",X"6D",X"DD",X"44",X"44",X"00",X"00",
		X"00",X"00",X"09",X"90",X"00",X"09",X"C6",X"69",X"99",X"99",X"99",X"C6",X"DD",X"66",X"66",X"66",
		X"DD",X"C4",X"50",X"00",X"00",X"00",X"00",X"0A",X"98",X"CD",X"89",X"90",X"00",X"00",X"00",X"00",
		X"6D",X"66",X"66",X"66",X"66",X"D8",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"99",X"88",X"89",
		X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"98",X"89",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"99",X"9A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A9",X"9A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"6A",X"00",X"00",X"00",X"00",X"00",X"E4",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"6D",X"65",X"E5",X"88",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"6D",X"D6",X"85",
		X"56",X"8D",X"DD",X"D8",X"90",X"0C",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"CD",X"DD",X"68",X"8E",X"88",X"DD",X"DD",X"DD",X"D8",X"00",X"6C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"66",X"C6",X"DD",X"D6",X"88",X"88",X"6C",X"88",X"89",X"99",X"6D",X"88",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"6D",X"C6",X"66",X"89",X"99",X"9D",X"D9",
		X"99",X"88",X"88",X"99",X"D6",X"DD",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"DD",X"D6",
		X"66",X"68",X"98",X"86",X"6F",X"F9",X"99",X"98",X"88",X"8D",X"DD",X"DD",X"DD",X"6C",X"00",X"00",
		X"00",X"4D",X"DD",X"DD",X"DD",X"DD",X"66",X"89",X"AC",X"C9",X"9F",X"FF",X"99",X"86",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"C0",X"00",X"56",X"66",X"6D",X"DD",X"DD",X"D6",X"68",X"96",X"CC",X"88",
		X"88",X"86",X"6D",X"D6",X"66",X"66",X"DD",X"DD",X"DD",X"D6",X"00",X"00",X"C6",X"66",X"66",X"6D",
		X"DD",X"D6",X"66",X"68",X"88",X"88",X"88",X"D6",X"66",X"DD",X"DD",X"66",X"DD",X"DD",X"DD",X"00",
		X"00",X"00",X"C6",X"66",X"66",X"66",X"DD",X"DD",X"88",X"82",X"28",X"88",X"C6",X"DD",X"DD",X"DD",
		X"D6",X"6D",X"DD",X"6C",X"00",X"00",X"0C",X"66",X"CC",X"C6",X"66",X"66",X"66",X"99",X"99",X"99",
		X"9C",X"6D",X"D6",X"66",X"6D",X"DD",X"55",X"5E",X"00",X"00",X"00",X"00",X"09",X"90",X"00",X"09",
		X"C6",X"69",X"99",X"99",X"99",X"C6",X"DD",X"66",X"66",X"66",X"DD",X"C5",X"E0",X"00",X"00",X"00",
		X"00",X"0A",X"98",X"CD",X"89",X"90",X"00",X"00",X"00",X"00",X"6D",X"66",X"66",X"66",X"66",X"D8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"99",X"88",X"89",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"98",X"89",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"99",X"9A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A9",X"9A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"11",X"11",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"FC",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"B0",X"00",X"CF",X"6F",X"60",X"6F",
		X"00",X"B0",X"00",X"00",X"00",X"0B",X"00",X"06",X"66",X"06",X"F6",X"FB",X"00",X"00",X"00",X"00",
		X"00",X"BC",X"F6",X"66",X"66",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"CF",X"66",X"66",X"66",
		X"60",X"60",X"00",X"00",X"00",X"00",X"0C",X"66",X"6B",X"66",X"66",X"66",X"00",X"00",X"00",X"00",
		X"00",X"00",X"CC",X"00",X"06",X"66",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",X"B6",
		X"6F",X"FC",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"66",X"00",X"6C",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"66",X"66",X"F6",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"66",X"FF",X"C0",
		X"0B",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"06",X"CC",X"00",X"0B",X"00",X"00",X"0B",X"00",
		X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",
		X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"0B",X"00",X"00",X"00",
		X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"F0",X"00",X"00",X"00",X"F6",X"00",X"00",X"00",X"00",X"00",X"06",
		X"60",X"00",X"00",X"06",X"F6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",
		X"60",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"60",X"00",X"0F",X"00",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"D0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"DD",
		X"F0",X"B0",X"00",X"00",X"00",X"00",X"06",X"66",X"60",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"6F",X"66",X"00",X"00",
		X"00",X"00",X"06",X"66",X"66",X"00",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"06",X"66",X"66",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"F0",X"00",X"00",X"06",X"00",
		X"60",X"00",X"D0",X"00",X"66",X"66",X"F0",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"06",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"0D",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"60",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"66",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"B0",X"00",X"00",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0B",X"00",X"0D",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"BB",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B0",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"D0",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D0",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"EE",X"EE",X"29",X"90",X"00",X"00",X"7E",X"EE",X"EE",
		X"29",X"90",X"00",X"00",X"7E",X"EE",X"EE",X"29",X"90",X"00",X"00",X"7E",X"EE",X"E2",X"29",X"90",
		X"00",X"00",X"CC",X"EE",X"CC",X"29",X"90",X"00",X"00",X"CC",X"CC",X"CC",X"C9",X"90",X"00",X"00",
		X"CC",X"CC",X"CC",X"C9",X"90",X"00",X"00",X"CC",X"CC",X"CC",X"C9",X"90",X"00",X"00",X"CC",X"CC",
		X"CC",X"C9",X"90",X"00",X"00",X"CC",X"CC",X"CC",X"C9",X"90",X"00",X"00",X"CC",X"CC",X"CC",X"C9",
		X"90",X"00",X"00",X"CC",X"CC",X"CC",X"29",X"90",X"00",X"00",X"7C",X"CC",X"CC",X"29",X"90",X"00",
		X"00",X"72",X"7C",X"C2",X"29",X"90",X"00",X"00",X"47",X"76",X"72",X"29",X"90",X"00",X"00",X"44",
		X"76",X"74",X"49",X"90",X"00",X"00",X"77",X"74",X"42",X"44",X"90",X"00",X"00",X"77",X"77",X"44",
		X"49",X"90",X"00",X"00",X"77",X"77",X"44",X"44",X"90",X"00",X"00",X"77",X"77",X"44",X"99",X"90",
		X"00",X"00",X"77",X"74",X"47",X"79",X"90",X"00",X"00",X"77",X"77",X"77",X"77",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"E2",X"29",X"90",X"00",X"00",X"EE",X"EE",X"EE",X"29",
		X"90",X"00",X"00",X"EE",X"EE",X"EE",X"29",X"90",X"00",X"00",X"EE",X"EE",X"EE",X"29",X"90",X"00",
		X"00",X"7E",X"EE",X"E2",X"29",X"90",X"00",X"00",X"7C",X"EE",X"22",X"29",X"90",X"00",X"00",X"7C",
		X"CC",X"C2",X"29",X"90",X"00",X"00",X"CC",X"CC",X"CC",X"29",X"90",X"00",X"00",X"CC",X"CC",X"CC",
		X"29",X"90",X"00",X"00",X"CC",X"CC",X"CC",X"C9",X"90",X"00",X"00",X"CC",X"CC",X"CC",X"C9",X"90",
		X"00",X"00",X"CC",X"CC",X"CC",X"C9",X"90",X"00",X"00",X"CC",X"CC",X"CC",X"CC",X"90",X"00",X"00",
		X"CC",X"CC",X"CC",X"CC",X"90",X"00",X"00",X"CC",X"CC",X"CC",X"CC",X"90",X"00",X"00",X"7C",X"CC",
		X"CC",X"C9",X"90",X"00",X"00",X"72",X"6C",X"CC",X"C9",X"90",X"00",X"00",X"26",X"92",X"2C",X"C9",
		X"90",X"00",X"00",X"47",X"99",X"96",X"29",X"90",X"00",X"00",X"44",X"79",X"99",X"69",X"90",X"00",
		X"00",X"77",X"47",X"79",X"69",X"90",X"00",X"00",X"77",X"77",X"44",X"29",X"90",X"00",X"00",X"00",
		X"00",X"04",X"44",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"40",X"00",X"00",X"00",X"00",X"00",
		X"40",X"40",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"28",X"43",X"29",X"20",X"31",X"39",
		X"38",X"34",X"2C",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",
		X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"00",X"09",X"92",
		X"EE",X"EE",X"E7",X"00",X"00",X"09",X"92",X"EE",X"EE",X"E7",X"00",X"00",X"09",X"92",X"EE",X"EE",
		X"E7",X"00",X"00",X"09",X"92",X"2E",X"EE",X"E7",X"00",X"00",X"09",X"92",X"CC",X"EE",X"CC",X"00",
		X"00",X"09",X"9C",X"CC",X"CC",X"CC",X"00",X"00",X"09",X"9C",X"CC",X"CC",X"CC",X"00",X"00",X"09",
		X"9C",X"CC",X"CC",X"CC",X"00",X"00",X"09",X"9C",X"CC",X"CC",X"CC",X"00",X"00",X"09",X"9C",X"CC",
		X"CC",X"CC",X"00",X"00",X"09",X"9C",X"CC",X"CC",X"CC",X"00",X"00",X"09",X"92",X"CC",X"CC",X"CC",
		X"00",X"00",X"09",X"92",X"CC",X"CC",X"C7",X"00",X"00",X"09",X"92",X"2C",X"C7",X"27",X"00",X"00",
		X"09",X"92",X"27",X"67",X"74",X"00",X"00",X"09",X"94",X"47",X"67",X"44",X"00",X"00",X"09",X"44",
		X"24",X"47",X"77",X"00",X"00",X"09",X"94",X"44",X"77",X"77",X"00",X"00",X"09",X"44",X"44",X"77",
		X"77",X"00",X"00",X"09",X"99",X"44",X"77",X"77",X"00",X"00",X"09",X"97",X"74",X"47",X"77",X"00",
		X"00",X"09",X"77",X"77",X"77",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"92",X"2E",
		X"EE",X"EE",X"00",X"00",X"09",X"92",X"EE",X"EE",X"EE",X"00",X"00",X"09",X"92",X"EE",X"EE",X"EE",
		X"00",X"00",X"09",X"92",X"EE",X"EE",X"EE",X"00",X"00",X"09",X"92",X"2E",X"EE",X"E0",X"00",X"00",
		X"09",X"92",X"22",X"EE",X"C0",X"00",X"00",X"09",X"92",X"2C",X"CC",X"C0",X"00",X"00",X"09",X"92",
		X"CC",X"CC",X"CC",X"00",X"00",X"09",X"92",X"CC",X"CC",X"CC",X"00",X"00",X"09",X"9C",X"CC",X"CC",
		X"CC",X"00",X"00",X"09",X"9C",X"CC",X"CC",X"CC",X"00",X"00",X"09",X"9C",X"CC",X"CC",X"CC",X"00",
		X"00",X"09",X"CC",X"CC",X"CC",X"CC",X"00",X"00",X"09",X"CC",X"CC",X"CC",X"CC",X"00",X"00",X"09",
		X"CC",X"CC",X"CC",X"CC",X"00",X"00",X"09",X"9C",X"CC",X"CC",X"C7",X"00",X"00",X"09",X"9C",X"CC",
		X"C6",X"27",X"00",X"00",X"09",X"9C",X"C2",X"29",X"62",X"00",X"00",X"09",X"92",X"69",X"99",X"74",
		X"00",X"00",X"09",X"96",X"99",X"97",X"44",X"00",X"00",X"09",X"96",X"97",X"74",X"77",X"00",X"00",
		X"09",X"92",X"44",X"77",X"77",X"00",X"00",X"00",X"44",X"40",X"00",X"00",X"00",X"00",X"04",X"40",
		X"40",X"00",X"00",X"00",X"00",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"EC",X"CC",X"E7",X"00",
		X"00",X"EC",X"CC",X"C7",X"00",X"00",X"EC",X"CC",X"C7",X"00",X"00",X"E2",X"CC",X"E7",X"00",X"00",
		X"EC",X"22",X"E7",X"00",X"00",X"CC",X"C2",X"E7",X"00",X"00",X"CC",X"CC",X"E7",X"00",X"0C",X"CC",
		X"CC",X"E7",X"00",X"0C",X"CC",X"CC",X"E7",X"00",X"0C",X"CC",X"CC",X"C7",X"00",X"0C",X"CC",X"CC",
		X"C7",X"00",X"0C",X"CC",X"CC",X"C7",X"00",X"04",X"EC",X"E7",X"C7",X"00",X"04",X"CE",X"77",X"47",
		X"00",X"00",X"40",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"E2",X"2E",X"77",X"00",
		X"00",X"E2",X"2E",X"7C",X"00",X"00",X"E2",X"2E",X"CC",X"00",X"00",X"E2",X"2E",X"CC",X"00",X"00",
		X"E2",X"AE",X"7C",X"00",X"00",X"EA",X"2E",X"CC",X"00",X"00",X"E2",X"2E",X"CC",X"00",X"00",X"E2",
		X"2E",X"CC",X"00",X"00",X"E2",X"2E",X"CC",X"00",X"00",X"E2",X"2E",X"CC",X"00",X"00",X"E2",X"2E",
		X"CC",X"00",X"00",X"E2",X"2E",X"CC",X"00",X"00",X"E2",X"EE",X"74",X"00",X"00",X"EE",X"77",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"92",X"22",X"27",
		X"77",X"00",X"00",X"09",X"92",X"22",X"27",X"77",X"00",X"00",X"09",X"92",X"22",X"2E",X"EE",X"00",
		X"00",X"09",X"92",X"22",X"EE",X"EE",X"00",X"00",X"09",X"92",X"22",X"EE",X"EE",X"00",X"00",X"09",
		X"92",X"22",X"EE",X"EE",X"00",X"00",X"09",X"92",X"2C",X"CE",X"EE",X"00",X"00",X"09",X"92",X"CC",
		X"CC",X"77",X"00",X"00",X"0F",X"9F",X"CC",X"CC",X"C7",X"00",X"0F",X"09",X"6C",X"6F",X"CC",X"CC",
		X"00",X"00",X"6C",X"EC",X"E6",X"CC",X"CC",X"00",X"F0",X"CE",X"CC",X"EC",X"FC",X"CC",X"00",X"06",
		X"CC",X"CC",X"C6",X"CC",X"CC",X"00",X"F0",X"EC",X"CC",X"EC",X"FC",X"C7",X"00",X"00",X"CC",X"CC",
		X"CC",X"CC",X"77",X"00",X"00",X"CC",X"CC",X"CC",X"CC",X"77",X"00",X"00",X"0C",X"CC",X"CC",X"CC",
		X"77",X"00",X"00",X"09",X"CC",X"CC",X"C7",X"77",X"00",X"00",X"09",X"9C",X"99",X"67",X"47",X"00",
		X"00",X"09",X"96",X"99",X"76",X"44",X"00",X"04",X"09",X"96",X"77",X"74",X"47",X"00",X"00",X"49",
		X"27",X"77",X"47",X"77",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"40",X"40",
		X"00",X"00",X"00",X"00",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"09",X"92",X"97",X"77",X"EE",
		X"00",X"00",X"09",X"92",X"97",X"77",X"EE",X"00",X"00",X"09",X"92",X"97",X"77",X"EE",X"00",X"00",
		X"09",X"92",X"97",X"77",X"EE",X"00",X"00",X"09",X"92",X"97",X"77",X"7E",X"00",X"00",X"09",X"92",
		X"97",X"77",X"7C",X"00",X"00",X"09",X"9C",X"C7",X"77",X"CC",X"00",X"00",X"09",X"9C",X"CC",X"C7",
		X"CC",X"00",X"00",X"09",X"92",X"CC",X"CF",X"CF",X"00",X"00",X"09",X"92",X"9F",X"CC",X"6C",X"00",
		X"00",X"09",X"92",X"97",X"6C",X"EC",X"00",X"00",X"09",X"92",X"F7",X"CE",X"CC",X"00",X"00",X"09",
		X"92",X"96",X"CC",X"CC",X"00",X"00",X"09",X"92",X"FC",X"EC",X"CC",X"00",X"00",X"09",X"92",X"9C",
		X"CC",X"CC",X"00",X"00",X"09",X"92",X"9C",X"CC",X"CC",X"00",X"00",X"09",X"92",X"77",X"CC",X"CC",
		X"00",X"00",X"09",X"99",X"77",X"76",X"CC",X"00",X"00",X"09",X"99",X"47",X"27",X"77",X"00",X"00",
		X"09",X"97",X"74",X"44",X"76",X"00",X"00",X"09",X"97",X"77",X"77",X"27",X"00",X"00",X"09",X"77",
		X"77",X"77",X"47",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"92",X"22",X"29",X"97",X"00",
		X"00",X"09",X"92",X"2C",X"29",X"97",X"00",X"00",X"09",X"92",X"22",X"C9",X"9C",X"00",X"00",X"09",
		X"92",X"2C",X"29",X"9C",X"00",X"00",X"09",X"92",X"C2",X"29",X"9C",X"00",X"00",X"09",X"92",X"22",
		X"99",X"9C",X"00",X"00",X"09",X"92",X"29",X"29",X"9C",X"00",X"00",X"09",X"92",X"92",X"C9",X"9C",
		X"00",X"00",X"09",X"99",X"22",X"C9",X"9C",X"00",X"00",X"09",X"92",X"2C",X"C9",X"9C",X"00",X"00",
		X"09",X"92",X"22",X"29",X"9C",X"00",X"00",X"09",X"92",X"2C",X"29",X"9C",X"00",X"00",X"09",X"92",
		X"22",X"C9",X"97",X"00",X"00",X"09",X"92",X"22",X"29",X"97",X"00",X"00",X"09",X"92",X"22",X"29",
		X"94",X"00",X"00",X"09",X"92",X"22",X"29",X"94",X"00",X"00",X"09",X"92",X"22",X"29",X"97",X"00",
		X"00",X"09",X"92",X"22",X"99",X"77",X"00",X"00",X"09",X"92",X"99",X"97",X"77",X"00",X"00",X"09",
		X"99",X"97",X"77",X"77",X"00",X"00",X"09",X"99",X"77",X"77",X"77",X"00",X"00",X"09",X"77",X"77",
		X"77",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"72",X"22",X"29",X"90",X"00",X"00",X"77",
		X"72",X"22",X"29",X"90",X"00",X"00",X"EE",X"E2",X"22",X"29",X"90",X"00",X"00",X"EE",X"EE",X"22",
		X"29",X"90",X"00",X"00",X"EE",X"EE",X"22",X"29",X"90",X"00",X"00",X"EE",X"EE",X"22",X"29",X"90",
		X"00",X"00",X"EE",X"EC",X"C2",X"29",X"90",X"00",X"00",X"77",X"CC",X"C2",X"29",X"90",X"00",X"00",
		X"7C",X"CC",X"CC",X"F9",X"F0",X"00",X"00",X"CC",X"CC",X"F6",X"C6",X"90",X"F0",X"00",X"CC",X"CC",
		X"6E",X"CE",X"C6",X"00",X"00",X"CC",X"CF",X"CE",X"CC",X"EC",X"0F",X"00",X"CC",X"CC",X"6C",X"CC",
		X"CE",X"60",X"00",X"7C",X"CF",X"CE",X"CC",X"CE",X"0F",X"00",X"77",X"CC",X"CC",X"CC",X"CC",X"00",
		X"00",X"77",X"CC",X"CC",X"CC",X"CC",X"00",X"00",X"77",X"CC",X"CC",X"CC",X"C0",X"00",X"00",X"77",
		X"7C",X"CC",X"CC",X"90",X"00",X"00",X"74",X"76",X"99",X"C9",X"90",X"00",X"00",X"44",X"67",X"99",
		X"69",X"90",X"00",X"00",X"74",X"47",X"77",X"69",X"90",X"40",X"00",X"77",X"74",X"77",X"72",X"94",
		X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"04",X"04",X"40",X"00",X"00",
		X"00",X"00",X"00",X"44",X"44",X"00",X"00",X"EE",X"77",X"79",X"29",X"90",X"00",X"00",X"EE",X"77",
		X"79",X"29",X"90",X"00",X"00",X"EE",X"77",X"79",X"29",X"90",X"00",X"00",X"EE",X"77",X"79",X"29",
		X"90",X"00",X"00",X"E7",X"77",X"79",X"29",X"90",X"00",X"00",X"C7",X"77",X"79",X"29",X"90",X"00",
		X"00",X"CC",X"77",X"7C",X"C9",X"90",X"00",X"00",X"CC",X"7C",X"CC",X"C9",X"90",X"00",X"00",X"FC",
		X"FC",X"CC",X"F9",X"90",X"00",X"00",X"C6",X"CC",X"F9",X"29",X"90",X"00",X"00",X"CE",X"C6",X"79",
		X"29",X"90",X"00",X"00",X"CC",X"EC",X"72",X"29",X"90",X"00",X"00",X"CC",X"CC",X"69",X"29",X"90",
		X"00",X"00",X"CC",X"CE",X"C2",X"29",X"90",X"00",X"00",X"CC",X"CC",X"C9",X"29",X"90",X"00",X"00",
		X"CC",X"CC",X"C9",X"29",X"90",X"00",X"00",X"CC",X"CC",X"77",X"29",X"90",X"00",X"00",X"CC",X"67",
		X"77",X"99",X"90",X"00",X"00",X"77",X"72",X"74",X"99",X"90",X"00",X"00",X"67",X"44",X"47",X"79",
		X"90",X"00",X"00",X"72",X"77",X"77",X"79",X"90",X"00",X"00",X"74",X"77",X"77",X"77",X"90",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"92",X"22",X"29",X"90",X"00",X"00",X"79",X"92",X"C2",
		X"29",X"90",X"00",X"00",X"C9",X"9C",X"22",X"29",X"90",X"00",X"00",X"C9",X"92",X"C2",X"29",X"90",
		X"00",X"00",X"C9",X"92",X"2C",X"29",X"90",X"00",X"00",X"C9",X"99",X"22",X"29",X"90",X"00",X"00",
		X"C9",X"92",X"92",X"29",X"90",X"00",X"00",X"C9",X"9C",X"29",X"29",X"90",X"00",X"00",X"C9",X"9C",
		X"22",X"99",X"90",X"00",X"00",X"C9",X"9C",X"C2",X"29",X"90",X"00",X"00",X"C9",X"92",X"22",X"29",
		X"90",X"00",X"00",X"C9",X"92",X"C2",X"29",X"90",X"00",X"00",X"79",X"9C",X"22",X"29",X"90",X"00",
		X"00",X"79",X"92",X"22",X"29",X"90",X"00",X"00",X"49",X"92",X"22",X"29",X"90",X"00",X"00",X"49",
		X"92",X"22",X"29",X"90",X"00",X"00",X"79",X"92",X"22",X"29",X"90",X"00",X"00",X"77",X"99",X"22",
		X"29",X"90",X"00",X"00",X"77",X"79",X"99",X"29",X"90",X"00",X"00",X"77",X"77",X"79",X"99",X"90",
		X"00",X"00",X"77",X"77",X"77",X"99",X"90",X"00",X"00",X"77",X"77",X"77",X"77",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"66",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"6A",
		X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"42",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"60",X"42",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"96",X"4B",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"66",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"00",X"99",X"66",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"06",
		X"90",X"9A",X"AA",X"00",X"96",X"00",X"00",X"00",X"00",X"00",X"06",X"9A",X"99",X"99",X"A9",X"96",
		X"60",X"00",X"00",X"00",X"00",X"68",X"A8",X"88",X"66",X"66",X"08",X"66",X"00",X"00",X"00",X"06",
		X"80",X"08",X"86",X"A6",X"66",X"00",X"86",X"60",X"00",X"0A",X"68",X"00",X"B8",X"86",X"66",X"66",
		X"B0",X"08",X"6A",X"00",X"06",X"80",X"0F",X"A8",X"86",X"A6",X"66",X"AF",X"00",X"68",X"00",X"06",
		X"80",X"BE",X"A8",X"66",X"66",X"66",X"AE",X"B0",X"68",X"00",X"06",X"80",X"FE",X"E0",X"66",X"A6",
		X"66",X"EE",X"F0",X"68",X"00",X"0A",X"A0",X"00",X"00",X"86",X"66",X"66",X"00",X"00",X"AA",X"00",
		X"CC",X"C0",X"00",X"00",X"98",X"99",X"90",X"00",X"0C",X"CC",X"00",X"C0",X"C0",X"00",X"00",X"0A",
		X"0A",X"00",X"00",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"0A",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CA",X"60",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"44",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"2A",X"3A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"04",X"2A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"04",
		X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"6B",X"B2",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"96",X"60",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"C9",
		X"96",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"99",X"AA",X"A9",X"C9",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"09",X"99",X"99",X"99",X"C6",X"C9",X"00",X"00",X"00",X"00",X"00",X"09",
		X"88",X"86",X"68",X"96",X"C0",X"00",X"00",X"00",X"00",X"00",X"C9",X"8A",X"66",X"68",X"96",X"60",
		X"00",X"00",X"00",X"00",X"00",X"C9",X"88",X"66",X"68",X"96",X"C6",X"F0",X"00",X"00",X"00",X"00",
		X"C9",X"8A",X"66",X"68",X"C9",X"C6",X"E0",X"00",X"00",X"00",X"00",X"6A",X"86",X"66",X"68",X"89",
		X"CC",X"0B",X"00",X"00",X"00",X"00",X"6A",X"9A",X"66",X"68",X"89",X"CC",X"EF",X"00",X"00",X"00",
		X"00",X"6A",X"98",X"66",X"88",X"89",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"89",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"A0",X"CC",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"A0",X"90",X"0C",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9C",X"C6",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"96",X"A6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C6",X"A6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"44",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"66",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"66",X"4A",X"3A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"04",
		X"2A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"04",X"22",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"6B",X"B2",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",
		X"96",X"60",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"96",X"60",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"6C",X"C9",X"AA",X"A9",X"98",X"00",X"00",X"00",X"00",X"00",X"09",X"6C",
		X"C9",X"99",X"9A",X"98",X"00",X"00",X"00",X"00",X"00",X"00",X"6C",X"98",X"86",X"66",X"DC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"6C",X"98",X"66",X"6A",X"DC",X"80",X"00",X"00",X"00",X"00",X"06",
		X"CC",X"98",X"66",X"66",X"DC",X"C0",X"00",X"00",X"00",X"00",X"B6",X"C9",X"C8",X"66",X"6A",X"D8",
		X"C0",X"00",X"00",X"00",X"0F",X"06",X"C9",X"C8",X"66",X"66",X"D8",X"C0",X"00",X"00",X"00",X"00",
		X"06",X"C9",X"86",X"66",X"6A",X"D8",X"C0",X"00",X"00",X"00",X"FE",X"EC",X"C9",X"98",X"66",X"66",
		X"D8",X"C0",X"00",X"00",X"00",X"00",X"00",X"AA",X"A9",X"89",X"99",X"A8",X"C0",X"00",X"00",X"00",
		X"00",X"0C",X"CC",X"00",X"A0",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"C0",X"00",X"A0",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"CC",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",
		X"0C",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0C",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"44",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"AA",X"06",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2B",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"2B",X"06",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"B6",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"29",X"66",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"00",X"99",X"66",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"06",X"90",X"9A",
		X"AA",X"00",X"96",X"00",X"00",X"00",X"00",X"00",X"06",X"9A",X"99",X"99",X"A9",X"96",X"60",X"00",
		X"00",X"00",X"00",X"68",X"A8",X"88",X"66",X"66",X"08",X"66",X"00",X"00",X"00",X"06",X"80",X"08",
		X"86",X"A6",X"66",X"00",X"86",X"60",X"00",X"0A",X"68",X"00",X"B8",X"86",X"66",X"66",X"B0",X"08",
		X"6A",X"00",X"06",X"80",X"0F",X"A8",X"86",X"A6",X"66",X"AF",X"00",X"68",X"00",X"06",X"80",X"BE",
		X"A8",X"66",X"66",X"66",X"AE",X"B0",X"68",X"00",X"06",X"80",X"FE",X"E0",X"66",X"A6",X"66",X"EE",
		X"F0",X"68",X"00",X"0A",X"A0",X"00",X"00",X"86",X"66",X"66",X"00",X"00",X"AA",X"00",X"CC",X"C0",
		X"00",X"00",X"98",X"99",X"90",X"00",X"0C",X"CC",X"00",X"C0",X"C0",X"00",X"00",X"0A",X"0A",X"00",
		X"00",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"0A",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"CC",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CA",X"60",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"44",X"44",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A3",X"03",X"66",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A2",X"BA",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"B0",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"2B",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"96",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"C9",X"96",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"99",X"AA",X"A9",X"C9",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"09",X"99",X"99",X"99",X"C6",X"C9",X"00",X"00",X"00",X"00",X"00",X"09",X"88",X"86",
		X"68",X"96",X"C0",X"00",X"00",X"00",X"00",X"00",X"C9",X"8A",X"66",X"68",X"96",X"60",X"00",X"00",
		X"00",X"00",X"00",X"C9",X"88",X"66",X"68",X"96",X"C6",X"F0",X"00",X"00",X"00",X"00",X"C9",X"8A",
		X"66",X"68",X"C9",X"C6",X"E0",X"00",X"00",X"00",X"00",X"6A",X"86",X"66",X"68",X"89",X"CC",X"0B",
		X"00",X"00",X"00",X"00",X"6A",X"9A",X"66",X"68",X"89",X"CC",X"EF",X"00",X"00",X"00",X"00",X"6A",
		X"98",X"66",X"88",X"89",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"89",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"A0",X"CC",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"90",X"0C",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9C",X"C6",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"96",X"A6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C6",X"A6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",
		X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A3",X"A3",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"BA",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"B0",X"66",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"2B",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"96",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"96",X"60",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"6C",X"C9",X"AA",X"A9",X"98",X"00",X"00",X"00",X"00",X"00",X"09",X"6C",X"C9",X"99",
		X"9A",X"98",X"00",X"00",X"00",X"00",X"00",X"00",X"6C",X"98",X"86",X"66",X"DC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"6C",X"98",X"66",X"6A",X"DC",X"80",X"00",X"00",X"00",X"00",X"06",X"CC",X"98",
		X"66",X"66",X"DC",X"C0",X"00",X"00",X"00",X"00",X"B6",X"C9",X"C8",X"66",X"6A",X"D8",X"C0",X"00",
		X"00",X"00",X"0F",X"06",X"C9",X"C8",X"66",X"66",X"D8",X"C0",X"00",X"00",X"00",X"00",X"06",X"C9",
		X"86",X"66",X"6A",X"D8",X"C0",X"00",X"00",X"00",X"FE",X"EC",X"C9",X"98",X"66",X"66",X"D8",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"AA",X"A9",X"89",X"99",X"A8",X"C0",X"00",X"00",X"00",X"00",X"0C",
		X"CC",X"00",X"A0",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"C0",X"00",X"A0",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"CC",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0C",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0C",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"44",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"44",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"AA",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"42",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"6A",
		X"42",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"AB",X"22",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"66",X"00",X"00",X"00",X"00",
		X"00",X"00",X"69",X"09",X"99",X"00",X"60",X"00",X"00",X"00",X"00",X"69",X"88",X"86",X"69",X"60",
		X"00",X"00",X"00",X"06",X"80",X"88",X"A6",X"60",X"86",X"00",X"00",X"00",X"68",X"0B",X"86",X"66",
		X"6B",X"08",X"60",X"00",X"06",X"80",X"FA",X"86",X"A6",X"60",X"F0",X"86",X"00",X"06",X"80",X"BA",
		X"C6",X"66",X"6A",X"B0",X"86",X"00",X"06",X"80",X"0A",X"C6",X"A6",X"6A",X"00",X"86",X"00",X"CC",
		X"C0",X"00",X"86",X"66",X"60",X"0C",X"CC",X"00",X"C0",X"C0",X"00",X"0A",X"0A",X"00",X"0C",X"0C",
		X"00",X"00",X"00",X"00",X"0A",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"66",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"44",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"33",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"42",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"6A",X"42",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"AB",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"69",X"68",X"C6",
		X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"98",X"C6",X"90",X"00",X"00",X"00",X"00",X"0C",X"66",
		X"66",X"98",X"60",X"00",X"00",X"00",X"00",X"0C",X"6A",X"66",X"98",X"60",X"00",X"00",X"00",X"00",
		X"0C",X"66",X"66",X"98",X"60",X"00",X"00",X"00",X"00",X"0C",X"6A",X"66",X"98",X"64",X"00",X"00",
		X"00",X"00",X"CC",X"66",X"66",X"98",X"6F",X"00",X"00",X"00",X"00",X"CC",X"9A",X"66",X"98",X"60",
		X"00",X"00",X"00",X"00",X"0C",X"99",X"89",X"CC",X"60",X"00",X"00",X"00",X"00",X"00",X"0A",X"0A",
		X"0C",X"60",X"00",X"00",X"00",X"00",X"00",X"0A",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"60",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"44",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"11",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"AA",X"42",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"6A",X"42",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"AB",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"CC",X"99",X"C0",X"00",X"00",X"00",X"00",X"00",X"8C",X"88",X"66",X"66",X"00",X"00",X"00",X"00",
		X"00",X"8C",X"86",X"6A",X"6D",X"00",X"00",X"00",X"00",X"00",X"8C",X"86",X"66",X"6D",X"00",X"00",
		X"00",X"00",X"04",X"8C",X"86",X"6A",X"6D",X"00",X"00",X"00",X"00",X"0B",X"8C",X"86",X"66",X"6D",
		X"00",X"00",X"00",X"00",X"00",X"8C",X"86",X"6A",X"6D",X"00",X"00",X"00",X"00",X"00",X"8C",X"86",
		X"89",X"6D",X"00",X"00",X"00",X"00",X"00",X"8C",X"0A",X"0A",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"C8",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"C8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"46",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"A6",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"A2",X"40",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"40",X"60",
		X"00",X"00",X"00",X"00",X"00",X"02",X"2B",X"A6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",
		X"69",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"69",X"00",X"00",X"00",X"00",X"00",X"00",
		X"69",X"09",X"99",X"00",X"60",X"00",X"00",X"00",X"00",X"69",X"88",X"86",X"69",X"60",X"00",X"00",
		X"00",X"06",X"80",X"88",X"A6",X"60",X"86",X"00",X"00",X"00",X"68",X"0B",X"86",X"66",X"6B",X"08",
		X"60",X"00",X"06",X"80",X"FA",X"86",X"A6",X"60",X"F0",X"86",X"00",X"06",X"80",X"BA",X"C6",X"66",
		X"6A",X"B0",X"86",X"00",X"06",X"80",X"0A",X"C6",X"A6",X"6A",X"00",X"86",X"00",X"CC",X"C0",X"00",
		X"86",X"66",X"60",X"0C",X"CC",X"00",X"C0",X"C0",X"00",X"0A",X"0A",X"00",X"0C",X"0C",X"00",X"00",
		X"00",X"00",X"0A",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"09",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"44",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"63",X"3A",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"A2",X"4A",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"4A",X"60",X"00",X"00",X"00",X"00",X"00",X"02",X"2B",X"A6",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"69",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"68",X"C6",X"00",X"00",
		X"00",X"00",X"00",X"09",X"99",X"98",X"C6",X"90",X"00",X"00",X"00",X"00",X"0C",X"66",X"66",X"98",
		X"60",X"00",X"00",X"00",X"00",X"0C",X"6A",X"66",X"98",X"60",X"00",X"00",X"00",X"00",X"0C",X"66",
		X"66",X"98",X"60",X"00",X"00",X"00",X"00",X"0C",X"6A",X"66",X"98",X"64",X"00",X"00",X"00",X"00",
		X"CC",X"66",X"66",X"98",X"6F",X"00",X"00",X"00",X"00",X"CC",X"9A",X"66",X"98",X"60",X"00",X"00",
		X"00",X"00",X"0C",X"99",X"89",X"CC",X"60",X"00",X"00",X"00",X"00",X"00",X"0A",X"0A",X"0C",X"60",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"60",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"44",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",
		X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"63",X"16",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"A2",X"4A",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"4A",X"60",X"00",X"00",X"00",
		X"00",X"00",X"02",X"2B",X"A6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"69",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"69",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"CC",X"99",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"8C",X"88",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"8C",
		X"86",X"6A",X"6D",X"00",X"00",X"00",X"00",X"00",X"8C",X"86",X"66",X"6D",X"00",X"00",X"00",X"00",
		X"04",X"8C",X"86",X"6A",X"6D",X"00",X"00",X"00",X"00",X"0B",X"8C",X"86",X"66",X"6D",X"00",X"00",
		X"00",X"00",X"00",X"8C",X"86",X"6A",X"6D",X"00",X"00",X"00",X"00",X"00",X"8C",X"86",X"89",X"6D",
		X"00",X"00",X"00",X"00",X"00",X"8C",X"0A",X"0A",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",
		X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"C8",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"C8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"46",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"40",X"00",X"00",X"00",X"00",X"00",X"06",
		X"66",X"00",X"00",X"00",X"00",X"00",X"66",X"AA",X"60",X"00",X"00",X"00",X"00",X"06",X"22",X"A0",
		X"00",X"00",X"00",X"00",X"06",X"AB",X"20",X"00",X"00",X"00",X"00",X"09",X"66",X"00",X"00",X"00",
		X"00",X"06",X"09",X"99",X"06",X"00",X"00",X"00",X"69",X"88",X"86",X"69",X"60",X"00",X"06",X"80",
		X"86",X"A6",X"60",X"86",X"00",X"68",X"0B",X"86",X"66",X"6B",X"08",X"60",X"68",X"0F",X"C6",X"A6",
		X"6F",X"08",X"60",X"6C",X"00",X"C6",X"66",X"60",X"0C",X"60",X"CC",X"00",X"86",X"66",X"60",X"0C",
		X"C0",X"00",X"00",X"0A",X"0A",X"00",X"00",X"00",X"00",X"00",X"0A",X"09",X"00",X"00",X"00",X"00",
		X"00",X"09",X"06",X"00",X"00",X"00",X"00",X"00",X"0C",X"06",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"66",X"60",X"00",X"00",X"00",X"00",X"C0",X"60",X"60",X"00",X"00",X"00",X"00",X"44",X"44",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"66",X"00",X"00",X"00",X"00",X"00",X"66",X"33",X"60",X"00",X"00",X"00",X"00",X"06",X"22",
		X"A0",X"00",X"00",X"00",X"00",X"06",X"AB",X"20",X"00",X"00",X"00",X"00",X"09",X"66",X"00",X"00",
		X"00",X"00",X"0C",X"C9",X"99",X"06",X"60",X"00",X"00",X"09",X"CC",X"C6",X"68",X"60",X"00",X"00",
		X"09",X"CA",X"66",X"69",X"60",X"00",X"00",X"09",X"C6",X"66",X"69",X"6B",X"00",X"00",X"09",X"CA",
		X"66",X"69",X"6F",X"00",X"00",X"09",X"C6",X"66",X"9C",X"C0",X"00",X"00",X"00",X"C6",X"66",X"9C",
		X"C0",X"00",X"00",X"00",X"0A",X"0A",X"00",X"00",X"00",X"00",X"00",X"0A",X"09",X"00",X"00",X"00",
		X"00",X"00",X"09",X"06",X"00",X"00",X"00",X"00",X"00",X"08",X"06",X"00",X"00",X"00",X"00",X"00",
		X"08",X"66",X"60",X"00",X"00",X"00",X"00",X"0C",X"60",X"60",X"00",X"00",X"00",X"00",X"CC",X"44",
		X"40",X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"44",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",X"00",X"00",X"00",
		X"00",X"66",X"33",X"60",X"00",X"00",X"00",X"00",X"06",X"22",X"A0",X"00",X"00",X"00",X"00",X"06",
		X"AB",X"20",X"00",X"00",X"00",X"00",X"09",X"66",X"00",X"00",X"00",X"00",X"06",X"09",X"99",X"C6",
		X"00",X"00",X"00",X"68",X"99",X"86",X"68",X"00",X"00",X"00",X"68",X"96",X"6A",X"68",X"00",X"00",
		X"0B",X"68",X"96",X"66",X"68",X"00",X"00",X"0F",X"68",X"96",X"6A",X"68",X"00",X"00",X"00",X"CC",
		X"96",X"66",X"68",X"00",X"00",X"00",X"CC",X"96",X"66",X"60",X"00",X"00",X"00",X"00",X"0A",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"09",X"00",X"00",X"00",X"00",X"00",X"09",X"08",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"C0",X"C8",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"C6",X"00",X"00",X"00",X"00",X"00",X"44",X"66",X"60",X"00",X"00",X"00",X"00",X"00",
		X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"44",X"40",X"00",X"00",X"00",X"00",X"06",X"66",X"00",
		X"00",X"00",X"00",X"00",X"6A",X"A6",X"60",X"00",X"00",X"00",X"00",X"02",X"2A",X"A0",X"00",X"00",
		X"00",X"00",X"2B",X"A6",X"00",X"00",X"00",X"00",X"00",X"06",X"69",X"00",X"00",X"00",X"00",X"06",
		X"09",X"99",X"06",X"00",X"00",X"00",X"69",X"88",X"86",X"69",X"60",X"00",X"06",X"80",X"86",X"A6",
		X"60",X"86",X"00",X"68",X"0B",X"86",X"66",X"6B",X"08",X"60",X"68",X"0F",X"C6",X"A6",X"6F",X"08",
		X"60",X"6C",X"00",X"C6",X"66",X"60",X"0C",X"60",X"CC",X"00",X"86",X"66",X"60",X"0C",X"C0",X"00",
		X"00",X"0A",X"0A",X"00",X"00",X"00",X"00",X"00",X"0A",X"09",X"00",X"00",X"00",X"00",X"00",X"09",
		X"06",X"00",X"00",X"00",X"00",X"00",X"0C",X"06",X"00",X"00",X"00",X"00",X"00",X"C0",X"66",X"60",
		X"00",X"00",X"00",X"00",X"C0",X"60",X"60",X"00",X"00",X"00",X"00",X"44",X"44",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",
		X"00",X"00",X"00",X"00",X"00",X"03",X"36",X"60",X"00",X"00",X"00",X"00",X"02",X"2A",X"A0",X"00",
		X"00",X"00",X"00",X"2B",X"A6",X"00",X"00",X"00",X"00",X"00",X"06",X"69",X"00",X"00",X"00",X"00",
		X"0C",X"C9",X"99",X"06",X"60",X"00",X"00",X"09",X"CC",X"C6",X"68",X"60",X"00",X"00",X"09",X"CA",
		X"66",X"69",X"60",X"00",X"00",X"09",X"C6",X"66",X"69",X"6B",X"00",X"00",X"09",X"CA",X"66",X"69",
		X"6F",X"00",X"00",X"09",X"C6",X"66",X"9C",X"C0",X"00",X"00",X"00",X"C6",X"66",X"9C",X"C0",X"00",
		X"00",X"00",X"0A",X"0A",X"00",X"00",X"00",X"00",X"00",X"0A",X"09",X"00",X"00",X"00",X"00",X"00",
		X"09",X"08",X"00",X"00",X"00",X"00",X"00",X"08",X"06",X"00",X"00",X"00",X"00",X"00",X"08",X"66",
		X"60",X"00",X"00",X"00",X"00",X"0C",X"60",X"60",X"00",X"00",X"00",X"00",X"C0",X"C4",X"40",X"00",
		X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"44",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",X"00",X"00",X"00",X"00",X"03",
		X"36",X"60",X"00",X"00",X"00",X"00",X"02",X"2A",X"A0",X"00",X"00",X"00",X"00",X"2B",X"A6",X"00",
		X"00",X"00",X"00",X"00",X"09",X"66",X"00",X"00",X"00",X"00",X"06",X"09",X"99",X"C6",X"00",X"00",
		X"00",X"68",X"99",X"86",X"68",X"00",X"00",X"00",X"68",X"96",X"6A",X"68",X"00",X"00",X"0B",X"68",
		X"96",X"66",X"68",X"00",X"00",X"0F",X"68",X"96",X"6A",X"68",X"00",X"00",X"00",X"CC",X"96",X"66",
		X"68",X"00",X"00",X"00",X"CC",X"96",X"66",X"60",X"00",X"00",X"00",X"00",X"0A",X"0A",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"09",X"00",X"00",X"00",X"00",X"00",X"09",X"08",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"C0",X"C8",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"C6",X"00",X"00",X"00",X"00",X"00",X"44",X"66",X"60",X"00",X"00",X"00",X"00",X"00",X"60",X"60",
		X"00",X"00",X"00",X"00",X"00",X"44",X"40",X"00",X"00",X"00",X"B0",X"00",X"0B",X"BB",X"00",X"BB",
		X"0B",X"B0",X"B0",X"00",X"B0",X"00",X"B0",X"00",X"0B",X"BB",X"00",X"BB",X"0B",X"B0",X"B0",X"00",
		X"B0",X"00",X"B0",X"00",X"0B",X"BB",X"00",X"BB",X"0B",X"B0",X"B0",X"00",X"B0",X"00",X"B0",X"00",
		X"0B",X"BB",X"00",X"BB",X"0B",X"B0",X"B0",X"00",X"B0",X"00",X"B0",X"00",X"0B",X"BB",X"00",X"BB",
		X"0B",X"B0",X"B0",X"00",X"B0",X"00",X"B0",X"00",X"0B",X"BB",X"00",X"BB",X"0B",X"B0",X"B0",X"00",
		X"B0",X"00",X"B0",X"00",X"0B",X"BB",X"00",X"BB",X"0B",X"B0",X"B0",X"00",X"B0",X"00",X"B0",X"00",
		X"0B",X"BB",X"00",X"BB",X"0B",X"B0",X"B0",X"00",X"B0",X"00",X"B0",X"00",X"0B",X"BB",X"00",X"BB",
		X"0B",X"B0",X"B0",X"00",X"B0",X"00",X"B0",X"00",X"0B",X"BB",X"00",X"BB",X"0B",X"B0",X"B0",X"00",
		X"B0",X"00",X"B0",X"00",X"0B",X"BB",X"00",X"BB",X"0B",X"B0",X"B0",X"00",X"B0",X"00",X"B0",X"00",
		X"0B",X"BB",X"00",X"BB",X"0B",X"B0",X"B0",X"00",X"B0",X"00",X"B0",X"00",X"0B",X"BB",X"00",X"BB",
		X"0B",X"B0",X"B0",X"00",X"B0",X"00",X"B0",X"00",X"0B",X"BB",X"00",X"BB",X"0B",X"B0",X"B0",X"00",
		X"B0",X"00",X"B0",X"00",X"0B",X"BB",X"00",X"BB",X"0B",X"B0",X"B0",X"00",X"B0",X"00",X"B0",X"00",
		X"0B",X"BB",X"00",X"BB",X"0B",X"B0",X"B0",X"00",X"B0",X"00",X"B0",X"00",X"0B",X"BB",X"00",X"BB",
		X"0B",X"B0",X"B0",X"00",X"B0",X"00",X"B0",X"00",X"0B",X"BB",X"00",X"BB",X"0B",X"B0",X"B0",X"00",
		X"B0",X"00",X"B0",X"00",X"0B",X"BB",X"00",X"BB",X"0B",X"B0",X"B0",X"00",X"B0",X"00",X"B0",X"00",
		X"0B",X"BB",X"00",X"BB",X"0B",X"B0",X"B0",X"00",X"B0",X"00",X"B0",X"00",X"0B",X"BB",X"00",X"BB",
		X"0B",X"B0",X"B0",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A9",X"88",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"88",X"99",
		X"90",X"98",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"98",X"99",X"99",X"48",X"89",X"94",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"89",X"99",X"99",X"89",X"99",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"98",X"99",X"99",X"98",X"99",
		X"99",X"94",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A9",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"89",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"90",
		X"09",X"89",X"99",X"98",X"00",X"00",X"98",X"88",X"99",X"99",X"99",X"94",X"00",X"0D",X"66",X"00",
		X"00",X"00",X"00",X"09",X"00",X"98",X"00",X"00",X"09",X"00",X"A9",X"88",X"89",X"99",X"99",X"99",
		X"99",X"00",X"88",X"C9",X"88",X"89",X"99",X"99",X"99",X"A9",X"80",X"00",X"00",X"99",X"98",X"88",
		X"88",X"88",X"88",X"88",X"88",X"99",X"00",X"88",X"9C",X"98",X"88",X"88",X"88",X"88",X"88",X"89",
		X"98",X"88",X"88",X"88",X"89",X"99",X"99",X"99",X"99",X"99",X"90",X"00",X"D9",X"98",X"88",X"89",
		X"99",X"99",X"98",X"88",X"99",X"99",X"CC",X"C9",X"99",X"99",X"98",X"88",X"88",X"88",X"88",X"88",
		X"00",X"DC",X"9D",X"88",X"98",X"88",X"88",X"99",X"98",X"88",X"99",X"AA",X"A9",X"9A",X"98",X"88",
		X"88",X"88",X"88",X"88",X"84",X"00",X"66",X"9D",X"89",X"88",X"88",X"88",X"88",X"99",X"98",X"89",
		X"99",X"99",X"A9",X"88",X"88",X"88",X"99",X"99",X"99",X"95",X"00",X"0C",X"66",X"98",X"88",X"99",
		X"98",X"88",X"89",X"99",X"99",X"99",X"9A",X"99",X"88",X"88",X"99",X"99",X"99",X"99",X"90",X"00",
		X"00",X"C6",X"68",X"89",X"AF",X"A9",X"98",X"88",X"99",X"99",X"99",X"9A",X"98",X"88",X"89",X"9A",
		X"AA",X"00",X"00",X"00",X"00",X"00",X"0C",X"C8",X"8A",X"AA",X"9A",X"A9",X"98",X"88",X"88",X"88",
		X"89",X"98",X"88",X"89",X"AA",X"99",X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"0A",X"9D",X"C9",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"98",X"DC",X"99",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"99",X"99",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"99",X"89",
		X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"A9",X"99",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A9",X"88",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"88",X"99",X"90",X"98",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"98",X"99",X"99",X"48",X"89",
		X"94",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"89",X"99",X"99",X"89",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"98",X"99",X"99",X"98",X"99",X"99",X"94",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"A9",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"89",X"99",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"90",X"09",X"89",X"99",X"98",X"00",X"00",X"98",
		X"88",X"99",X"99",X"99",X"94",X"00",X"0D",X"66",X"00",X"00",X"00",X"00",X"09",X"00",X"98",X"00",
		X"00",X"09",X"00",X"A9",X"88",X"89",X"99",X"99",X"99",X"99",X"00",X"88",X"C9",X"88",X"89",X"99",
		X"99",X"99",X"A9",X"80",X"00",X"00",X"99",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"99",X"00",
		X"88",X"9C",X"98",X"88",X"88",X"88",X"88",X"88",X"89",X"98",X"88",X"88",X"88",X"89",X"99",X"99",
		X"99",X"99",X"99",X"90",X"00",X"D9",X"98",X"88",X"89",X"99",X"99",X"98",X"88",X"99",X"99",X"CC",
		X"C9",X"99",X"99",X"98",X"88",X"88",X"88",X"88",X"88",X"00",X"DC",X"9D",X"88",X"98",X"88",X"88",
		X"99",X"98",X"88",X"99",X"AA",X"A9",X"9A",X"98",X"88",X"88",X"88",X"88",X"88",X"84",X"00",X"66",
		X"9D",X"89",X"88",X"88",X"88",X"88",X"99",X"98",X"89",X"99",X"99",X"A9",X"88",X"88",X"88",X"99",
		X"99",X"99",X"95",X"00",X"0C",X"66",X"98",X"88",X"99",X"98",X"88",X"89",X"99",X"99",X"99",X"9A",
		X"99",X"88",X"88",X"99",X"99",X"99",X"99",X"90",X"00",X"00",X"C6",X"68",X"89",X"AA",X"A9",X"98",
		X"88",X"99",X"99",X"99",X"9A",X"98",X"88",X"89",X"9A",X"AA",X"99",X"A0",X"00",X"00",X"00",X"0C",
		X"C8",X"8A",X"9D",X"C9",X"99",X"98",X"88",X"88",X"88",X"89",X"98",X"88",X"8A",X"98",X"DC",X"99",
		X"A0",X"00",X"00",X"00",X"00",X"00",X"0A",X"99",X"99",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"99",X"89",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A9",X"99",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"88",X"9A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"89",X"09",X"99",X"88",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"49",X"98",X"84",X"99",
		X"99",X"89",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"98",X"99",X"99",X"98",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"49",X"99",X"99",X"89",X"99",X"99",X"89",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"99",X"98",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"9A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"49",X"99",X"99",X"99",X"88",X"89",X"00",X"00",X"89",X"99",X"98",X"90",X"09",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"99",X"99",X"98",X"88",X"9A",X"00",X"90",X"00",X"00",
		X"89",X"00",X"90",X"00",X"00",X"00",X"00",X"66",X"D0",X"00",X"99",X"88",X"88",X"88",X"88",X"88",
		X"88",X"89",X"99",X"00",X"00",X"08",X"9A",X"99",X"99",X"99",X"98",X"88",X"9C",X"88",X"00",X"09",
		X"99",X"99",X"99",X"99",X"99",X"98",X"88",X"88",X"88",X"89",X"98",X"88",X"88",X"88",X"88",X"88",
		X"89",X"C9",X"88",X"00",X"88",X"88",X"88",X"88",X"88",X"89",X"99",X"99",X"9C",X"CC",X"99",X"99",
		X"88",X"89",X"99",X"99",X"98",X"88",X"89",X"9D",X"00",X"48",X"88",X"88",X"88",X"88",X"88",X"89",
		X"A9",X"9A",X"AA",X"99",X"88",X"89",X"99",X"88",X"88",X"89",X"88",X"D9",X"CD",X"00",X"59",X"99",
		X"99",X"99",X"88",X"88",X"88",X"9A",X"99",X"99",X"98",X"89",X"99",X"88",X"88",X"88",X"88",X"98",
		X"D9",X"66",X"00",X"09",X"99",X"99",X"99",X"99",X"88",X"88",X"99",X"A9",X"99",X"99",X"99",X"98",
		X"88",X"89",X"99",X"88",X"89",X"66",X"C0",X"00",X"00",X"00",X"00",X"AA",X"A9",X"98",X"88",X"89",
		X"A9",X"99",X"99",X"99",X"88",X"89",X"9A",X"FA",X"98",X"86",X"6C",X"00",X"00",X"00",X"0A",X"AA",
		X"99",X"AA",X"98",X"88",X"89",X"98",X"88",X"88",X"88",X"89",X"9A",X"A9",X"AA",X"A8",X"8C",X"C0",
		X"00",X"00",X"00",X"0A",X"99",X"CD",X"89",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",
		X"9C",X"D9",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"98",X"99",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"99",X"99",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"99",
		X"9A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"88",X"9A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"89",X"09",X"99",X"88",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"49",X"98",X"84",X"99",X"99",X"89",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"98",X"99",X"99",X"98",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"49",
		X"99",X"99",X"89",X"99",X"99",X"89",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"99",X"99",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"9A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"49",X"99",X"99",X"99",X"88",X"89",X"00",
		X"00",X"89",X"99",X"98",X"90",X"09",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",
		X"99",X"99",X"98",X"88",X"9A",X"00",X"90",X"00",X"00",X"89",X"00",X"90",X"00",X"00",X"00",X"00",
		X"66",X"D0",X"00",X"99",X"88",X"88",X"88",X"88",X"88",X"88",X"89",X"99",X"00",X"00",X"08",X"9A",
		X"99",X"99",X"99",X"98",X"88",X"9C",X"88",X"00",X"09",X"99",X"99",X"99",X"99",X"99",X"98",X"88",
		X"88",X"88",X"89",X"98",X"88",X"88",X"88",X"88",X"88",X"89",X"C9",X"88",X"00",X"88",X"88",X"88",
		X"88",X"88",X"89",X"99",X"99",X"9C",X"CC",X"99",X"99",X"88",X"89",X"99",X"99",X"98",X"88",X"89",
		X"9D",X"00",X"48",X"88",X"88",X"88",X"88",X"88",X"89",X"A9",X"9A",X"AA",X"99",X"88",X"89",X"99",
		X"88",X"88",X"89",X"88",X"D9",X"CD",X"00",X"59",X"99",X"99",X"99",X"88",X"88",X"88",X"9A",X"99",
		X"99",X"98",X"89",X"99",X"88",X"88",X"88",X"88",X"98",X"D9",X"66",X"00",X"09",X"99",X"99",X"99",
		X"99",X"88",X"88",X"99",X"A9",X"99",X"99",X"99",X"98",X"88",X"89",X"99",X"88",X"89",X"66",X"C0",
		X"00",X"00",X"0A",X"99",X"AA",X"A9",X"98",X"88",X"89",X"A9",X"99",X"99",X"99",X"88",X"89",X"9A",
		X"AA",X"98",X"86",X"6C",X"00",X"00",X"00",X"0A",X"99",X"CD",X"89",X"A8",X"88",X"89",X"98",X"88",
		X"88",X"88",X"89",X"99",X"9C",X"D9",X"A8",X"8C",X"C0",X"00",X"00",X"00",X"00",X"99",X"98",X"99",
		X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"99",X"99",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"99",X"9A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"CC",X"E0",X"00",X"00",X"00",X"CC",
		X"E0",X"00",X"00",X"00",X"CC",X"E0",X"00",X"00",X"00",X"CC",X"CE",X"00",X"00",X"00",X"00",X"CE",
		X"00",X"00",X"00",X"0C",X"CC",X"E0",X"00",X"00",X"0C",X"CC",X"CE",X"00",X"00",X"CC",X"CC",X"CC",
		X"F0",X"00",X"CC",X"CC",X"CC",X"EF",X"00",X"CC",X"CC",X"CC",X"E6",X"00",X"CC",X"CC",X"CC",X"E6",
		X"00",X"CC",X"CC",X"CC",X"CF",X"00",X"CC",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"CC",X"00",X"00",
		X"CC",X"CC",X"E0",X"00",X"00",X"C0",X"EE",X"00",X"00",X"00",X"C0",X"0C",X"C0",X"00",X"00",X"00",
		X"00",X"C0",X"C0",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"0C",X"CC",X"00",X"00",X"00",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"0E",X"CC",X"00",X"00",X"00",X"0E",
		X"CC",X"00",X"00",X"00",X"0E",X"CC",X"00",X"00",X"00",X"EC",X"CC",X"00",X"00",X"00",X"EC",X"00",
		X"00",X"00",X"0E",X"CC",X"C0",X"00",X"00",X"EC",X"CC",X"C0",X"00",X"0F",X"CC",X"CC",X"CC",X"00",
		X"FE",X"CC",X"CC",X"CC",X"00",X"6E",X"CC",X"CC",X"CC",X"00",X"6E",X"CC",X"CC",X"CC",X"00",X"FC",
		X"CC",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"CC",X"00",X"00",X"0E",
		X"CC",X"CC",X"00",X"00",X"00",X"EE",X"0C",X"00",X"00",X"0C",X"C0",X"0C",X"00",X"0C",X"0C",X"00",
		X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"CC",X"C0",X"00",X"00",X"00",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"C8",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"99",X"99",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"97",X"79",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"AA",X"A4",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"B5",X"AA",X"A7",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"05",X"A7",X"77",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"07",X"74",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"77",X"75",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"EE",
		X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"55",X"55",X"50",X"00",X"00",
		X"00",X"00",X"0C",X"00",X"00",X"CA",X"0E",X"55",X"E0",X"5E",X"00",X"00",X"00",X"00",X"CC",X"CC",
		X"CC",X"C5",X"5E",X"E5",X"E0",X"05",X"00",X"00",X"00",X"00",X"99",X"99",X"EE",X"CC",X"E5",X"55",
		X"E0",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"94",X"EE",X"54",X"5E",X"E0",X"5E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"EA",X"5E",X"E4",X"55",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"E5",X"E4",X"5E",X"05",X"0E",X"E5",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"E5",
		X"E0",X"00",X"0E",X"0E",X"E0",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"45",X"00",X"00",X"0E",
		X"50",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"0B",X"50",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"E0",X"00",X"00",X"BB",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"B4",X"00",X"00",
		X"00",X"0E",X"BB",X"B5",X"00",X"00",X"00",X"00",X"0B",X"00",X"40",X"00",X"00",X"00",X"00",X"5B",
		X"B0",X"00",X"00",X"0B",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",
		X"00",X"00",X"98",X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"8C",
		X"89",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"89",X"99",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"77",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EA",X"AA",X"47",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2B",X"5A",X"AA",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"5A",X"77",X"70",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"07",X"75",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"75",
		X"5E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"EE",X"54",X"50",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"55",X"5E",X"55",X"00",X"00",X"00",X"0C",X"00",X"00",
		X"CA",X"00",X"0E",X"55",X"5E",X"05",X"E0",X"00",X"00",X"CC",X"CC",X"CC",X"C5",X"5E",X"AE",X"E5",
		X"E0",X"00",X"50",X"00",X"00",X"99",X"99",X"EE",X"CC",X"8A",X"E5",X"55",X"E0",X"00",X"50",X"00",
		X"00",X"00",X"09",X"C4",X"EE",X"9A",X"54",X"55",X"EE",X"E5",X"E0",X"0E",X"00",X"00",X"00",X"05",
		X"EC",X"9A",X"55",X"5E",X"E4",X"EE",X"00",X"E5",X"E0",X"00",X"00",X"00",X"CC",X"90",X"E5",X"5E",
		X"E4",X"5E",X"0E",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"0E",X"E5",X"AE",X"E0",X"00",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E4",X"40",X"00",X"0E",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"B4",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5B",X"BB",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"88",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"C8",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"99",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"97",X"79",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"AA",X"A4",X"70",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"B5",X"AA",X"A7",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",
		X"05",X"A7",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"07",X"74",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"77",X"75",X"5E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"EE",X"54",X"5E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"05",X"55",X"5E",X"55",X"50",X"00",X"00",X"0C",X"00",X"00",X"CA",X"00",X"0E",X"55",
		X"5E",X"00",X"55",X"00",X"00",X"CC",X"CC",X"CC",X"C5",X"5E",X"AE",X"E5",X"E0",X"00",X"05",X"00",
		X"00",X"99",X"99",X"EE",X"CC",X"8A",X"E5",X"55",X"E0",X"0E",X"E5",X"00",X"00",X"00",X"09",X"C4",
		X"EE",X"9A",X"54",X"55",X"50",X"E4",X"EE",X"00",X"00",X"00",X"00",X"05",X"EC",X"9A",X"55",X"55",
		X"55",X"E4",X"5E",X"0E",X"00",X"00",X"00",X"00",X"CC",X"90",X"E5",X"55",X"EE",X"AE",X"E0",X"E5",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"0E",X"E5",X"4E",X"E0",X"00",X"00",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"BB",X"40",X"00",X"00",X"0E",X"50",X"00",X"00",X"00",X"00",X"00",X"0B",X"B0",
		X"E5",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"0E",X"50",X"0E",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"E5",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"4B",X"B0",X"00",X"05",X"55",X"00",X"00",X"00",X"00",X"00",X"0B",X"5B",X"B5",X"00",
		X"E5",X"5E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"88",X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"A2",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"BB",X"BE",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"7B",X"75",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E7",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"45",X"E4",X"E5",X"4E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"E5",X"5E",X"55",
		X"E5",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"5E",X"CE",X"E5",X"55",X"00",X"5E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"5C",X"6C",X"E5",X"5E",X"00",X"0E",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"58",X"A8",X"E4",X"55",X"EE",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"89",X"AE",X"45",
		X"5E",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"EE",X"A5",X"55",X"50",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"5E",X"E5",X"55",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"5E",X"5E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"B0",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"B4",X"B5",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"5B",X"50",X"5B",X"5B",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"88",X"89",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"98",X"C8",X"88",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"98",X"88",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"77",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"74",X"AA",X"AE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"AA",
		X"A5",X"B2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"77",X"A5",X"0B",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"E4",X"77",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"55",X"77",X"70",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"4E",X"E5",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"50",X"E5",X"5E",X"0A",X"C0",X"00",X"0C",X"00",X"00",X"00",X"00",X"05",
		X"00",X"E5",X"EE",X"55",X"CC",X"CC",X"CC",X"C0",X"00",X"00",X"00",X"05",X"00",X"E5",X"55",X"EC",
		X"CE",X"E9",X"99",X"90",X"00",X"00",X"00",X"0E",X"50",X"EE",X"54",X"5E",X"E4",X"C9",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E5",X"54",X"EE",X"5C",X"E5",X"00",X"00",X"00",X"00",X"05",X"EE",X"05",
		X"0E",X"54",X"E5",X"EC",X"C0",X"00",X"00",X"00",X"00",X"EE",X"0E",X"00",X"00",X"E5",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"5E",X"00",X"00",X"05",X"40",X"05",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"5B",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"0B",
		X"B0",X"00",X"00",X"E4",X"00",X"00",X"00",X"00",X"00",X"05",X"BB",X"BE",X"00",X"00",X"00",X"04",
		X"B0",X"00",X"00",X"00",X"00",X"BB",X"50",X"00",X"00",X"00",X"00",X"40",X"0B",X"00",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4B",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"88",X"88",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"8C",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"99",X"88",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"97",X"79",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"4A",X"AA",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"7A",X"AA",
		X"5B",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"7A",X"50",X"B0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"70",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"77",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"55",X"7E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"5E",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"05",X"5E",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E5",
		X"0E",X"55",X"5E",X"00",X"0A",X"C0",X"00",X"0C",X"00",X"00",X"00",X"50",X"00",X"E5",X"EE",X"AE",
		X"55",X"CC",X"CC",X"CC",X"C0",X"00",X"00",X"50",X"00",X"E5",X"55",X"EA",X"8C",X"CE",X"E9",X"99",
		X"90",X"0E",X"00",X"E5",X"EE",X"E5",X"54",X"5A",X"9E",X"E4",X"C9",X"00",X"00",X"E5",X"E0",X"0E",
		X"E4",X"EE",X"55",X"5A",X"9C",X"E5",X"00",X"00",X"00",X"50",X"0E",X"0E",X"54",X"EE",X"55",X"E0",
		X"9C",X"C0",X"00",X"00",X"00",X"0E",X"00",X"00",X"EE",X"A5",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"44",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"E0",X"00",
		X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"B5",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"4B",X"BB",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"89",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"98",X"C8",X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"98",X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"77",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"74",X"AA",X"AE",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"AA",X"A5",X"B2",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"77",X"A5",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"E4",X"77",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"55",X"77",X"70",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"54",X"5E",X"E5",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",
		X"5E",X"55",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"50",X"0E",X"55",X"5E",X"00",
		X"0A",X"C0",X"00",X"0C",X"00",X"00",X"05",X"00",X"00",X"E5",X"EE",X"AE",X"55",X"CC",X"CC",X"CC",
		X"C0",X"00",X"05",X"EE",X"00",X"E5",X"55",X"EA",X"8C",X"CE",X"E9",X"99",X"90",X"00",X"0E",X"E4",
		X"E0",X"55",X"54",X"5A",X"9E",X"E4",X"C9",X"00",X"00",X"0E",X"0E",X"54",X"E5",X"55",X"55",X"5A",
		X"9C",X"E5",X"00",X"00",X"00",X"E5",X"E0",X"EE",X"AE",X"E5",X"55",X"E0",X"9C",X"C0",X"00",X"00",
		X"00",X"E0",X"00",X"00",X"EE",X"45",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"5E",X"00",X"00",
		X"00",X"4B",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"05",X"E0",X"BB",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"5E",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"05",X"E0",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"55",
		X"00",X"00",X"BB",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"55",X"E0",X"05",X"BB",
		X"5B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"C9",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"89",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"A4",X"79",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"5A",X"A7",X"70",X"00",X"00",X"00",
		X"00",X"00",X"00",X"B0",X"57",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"7E",
		X"E5",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"57",X"75",X"4E",X"00",X"00",X"00",X"00",
		X"0C",X"00",X"0C",X"05",X"5E",X"55",X"00",X"00",X"00",X"00",X"CC",X"CC",X"CC",X"55",X"55",X"05",
		X"00",X"00",X"00",X"00",X"99",X"99",X"5C",X"EE",X"5E",X"05",X"E0",X"00",X"00",X"00",X"00",X"09",
		X"4E",X"54",X"55",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"5E",X"E4",X"45",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"5E",X"E5",X"5A",X"EE",X"5E",X"00",X"00",X"00",X"00",X"00",X"0E",
		X"EE",X"00",X"0E",X"0E",X"E0",X"00",X"00",X"00",X"00",X"50",X"4B",X"00",X"00",X"0E",X"50",X"00",
		X"00",X"00",X"04",X"00",X"05",X"B5",X"0B",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"0B",
		X"BB",X"B5",X"00",X"00",X"00",X"0B",X"04",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"0B",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"98",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"88",X"8C",X"90",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"99",
		X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"AA",X"47",X"90",X"00",X"00",X"00",X"00",
		X"00",X"0B",X"B5",X"AA",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"05",X"77",X"70",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"07",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"75",X"4E",X"00",X"00",
		X"00",X"0C",X"00",X"0C",X"00",X"05",X"55",X"55",X"E0",X"00",X"00",X"CC",X"CC",X"CC",X"5E",X"05",
		X"55",X"0E",X"50",X"00",X"00",X"99",X"99",X"5C",X"CA",X"EE",X"50",X"00",X"5E",X"00",X"00",X"00",
		X"09",X"45",X"9E",X"54",X"55",X"00",X"50",X"00",X"00",X"00",X"00",X"55",X"9E",X"55",X"5E",X"44",
		X"50",X"E0",X"00",X"00",X"00",X"0C",X"9E",X"55",X"5A",X"55",X"0E",X"5E",X"00",X"00",X"00",X"00",
		X"00",X"E4",X"5E",X"E0",X"0E",X"0E",X"50",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"BB",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"BB",X"B5",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"89",X"99",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"AA",X"A4",X"79",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"5A",X"A7",
		X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"57",X"77",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"7E",X"E5",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"57",X"75",X"45",
		X"00",X"00",X"00",X"0C",X"00",X"0C",X"00",X"05",X"55",X"0E",X"50",X"00",X"00",X"CC",X"CC",X"CC",
		X"5E",X"05",X"55",X"00",X"E5",X"00",X"00",X"99",X"99",X"5C",X"CA",X"EE",X"5E",X"00",X"05",X"00",
		X"00",X"00",X"09",X"45",X"9E",X"54",X"55",X"04",X"4E",X"05",X"00",X"00",X"00",X"55",X"9E",X"55",
		X"5A",X"E5",X"50",X"00",X"E0",X"00",X"00",X"0C",X"9E",X"55",X"5E",X"E0",X"00",X"EE",X"50",X"00",
		X"00",X"00",X"00",X"E4",X"B4",X"00",X"0E",X"E0",X"00",X"00",X"00",X"00",X"00",X"B4",X"E5",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"50",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"B0",X"00",X"00",X"55",X"00",
		X"00",X"00",X"00",X"B5",X"BB",X"E0",X"05",X"55",X"E0",X"00",X"00",X"00",X"00",X"00",X"0A",X"88",
		X"8A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"52",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"7B",X"74",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E7",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"47",
		X"45",X"50",X"00",X"00",X"00",X"00",X"00",X"05",X"C0",X"5E",X"5E",X"E5",X"00",X"00",X"00",X"00",
		X"00",X"59",X"C9",X"E5",X"50",X"00",X"50",X"00",X"00",X"00",X"00",X"5C",X"A8",X"E5",X"5E",X"00",
		X"E5",X"00",X"00",X"00",X"00",X"09",X"89",X"E4",X"45",X"E5",X"40",X"00",X"00",X"00",X"00",X"05",
		X"AE",X"E5",X"45",X"AE",X"50",X"00",X"00",X"00",X"00",X"00",X"E5",X"55",X"55",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"5E",X"5E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"B0",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B4",X"B0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"B5",X"B0",X"B5",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"89",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"C8",X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"99",
		X"99",X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"09",X"74",X"AA",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"77",X"AA",X"5B",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"77",X"50",
		X"B0",X"00",X"00",X"00",X"00",X"00",X"E5",X"EE",X"70",X"40",X"00",X"00",X"00",X"00",X"00",X"0E",
		X"45",X"77",X"50",X"40",X"00",X"00",X"00",X"00",X"00",X"05",X"5E",X"55",X"0C",X"00",X"0C",X"00",
		X"00",X"00",X"00",X"05",X"05",X"55",X"5C",X"CC",X"CC",X"C0",X"00",X"00",X"00",X"E5",X"0E",X"5E",
		X"EC",X"59",X"99",X"90",X"00",X"00",X"00",X"05",X"05",X"54",X"5E",X"49",X"00",X"00",X"00",X"00",
		X"00",X"05",X"44",X"EE",X"5E",X"50",X"00",X"00",X"00",X"0E",X"5E",X"EA",X"55",X"EE",X"5E",X"00",
		X"00",X"00",X"00",X"EE",X"0E",X"00",X"0E",X"EE",X"00",X"00",X"00",X"00",X"00",X"5E",X"00",X"00",
		X"0B",X"40",X"50",X"00",X"00",X"00",X"00",X"00",X"0B",X"05",X"B5",X"00",X"04",X"00",X"00",X"00",
		X"00",X"05",X"BB",X"BB",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",
		X"04",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4B",X"00",X"00",X"00",
		X"00",X"00",X"08",X"88",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9C",X"88",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"98",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"97",X"4A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"7A",X"A5",X"BB",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"77",X"75",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"57",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"45",X"75",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E5",X"55",X"55",X"00",X"0C",
		X"00",X"0C",X"00",X"00",X"00",X"5E",X"05",X"55",X"0E",X"5C",X"CC",X"CC",X"C0",X"00",X"0E",X"50",
		X"00",X"5E",X"EA",X"CC",X"59",X"99",X"90",X"00",X"00",X"50",X"05",X"54",X"5E",X"95",X"49",X"00",
		X"00",X"00",X"E0",X"54",X"4E",X"55",X"5E",X"95",X"50",X"00",X"00",X"0E",X"5E",X"05",X"5A",X"55",
		X"5E",X"9C",X"00",X"00",X"00",X"5E",X"0E",X"00",X"EE",X"54",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5B",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"4B",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",
		X"BB",X"B5",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",
		X"89",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"C8",X"88",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"99",X"99",X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"09",X"74",X"AA",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"AA",X"5B",X"B0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"77",X"50",X"B0",X"00",X"00",X"00",X"00",X"00",X"E5",X"EE",X"70",X"40",X"00",X"00",
		X"00",X"00",X"00",X"05",X"45",X"77",X"50",X"40",X"00",X"00",X"00",X"00",X"00",X"5E",X"05",X"55",
		X"00",X"0C",X"00",X"0C",X"00",X"00",X"05",X"E0",X"05",X"55",X"0E",X"5C",X"CC",X"CC",X"C0",X"00",
		X"05",X"00",X"0E",X"5E",X"EA",X"CC",X"59",X"99",X"90",X"05",X"0E",X"44",X"05",X"54",X"5E",X"95",
		X"49",X"00",X"00",X"E0",X"00",X"55",X"EA",X"55",X"5E",X"95",X"50",X"00",X"00",X"5E",X"E0",X"00",
		X"EE",X"55",X"5E",X"9C",X"00",X"00",X"00",X"00",X"EE",X"00",X"04",X"B4",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E5",X"E4",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",
		X"5B",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",
		X"05",X"50",X"00",X"00",X"B4",X"00",X"00",X"00",X"00",X"00",X"00",X"E5",X"55",X"00",X"EB",X"B5",
		X"B0",X"00",X"00",X"00",X"00",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"FF",X"98",X"88",
		X"8F",X"00",X"00",X"00",X"00",X"0F",X"88",X"89",X"99",X"8F",X"00",X"00",X"00",X"00",X"0F",X"FF",
		X"AA",X"77",X"F0",X"00",X"00",X"00",X"00",X"FE",X"BE",X"AA",X"77",X"F0",X"00",X"00",X"00",X"00",
		X"0F",X"F5",X"77",X"4F",X"FF",X"00",X"00",X"00",X"00",X"00",X"F4",X"F7",X"FF",X"5E",X"F0",X"00",
		X"00",X"00",X"00",X"0F",X"0F",X"77",X"54",X"5F",X"00",X"00",X"00",X"00",X"FF",X"FC",X"F5",X"5F",
		X"E5",X"F0",X"00",X"00",X"0F",X"CC",X"CC",X"5E",X"5E",X"F5",X"F0",X"00",X"00",X"0F",X"99",X"95",
		X"E4",X"EE",X"5E",X"F0",X"00",X"00",X"00",X"FF",X"F4",X"5E",X"54",X"EF",X"00",X"00",X"00",X"00",
		X"00",X"FE",X"EA",X"5E",X"AE",X"E5",X"00",X"00",X"00",X"00",X"0F",X"5E",X"4F",X"F0",X"E0",X"50",
		X"00",X"00",X"00",X"F5",X"FF",X"FB",X"FF",X"00",X"00",X"00",X"00",X"0F",X"4F",X"00",X"0F",X"4B",
		X"FF",X"00",X"00",X"00",X"F4",X"E4",X"00",X"00",X"FF",X"B5",X"F0",X"00",X"00",X"BF",X"FF",X"00",
		X"00",X"00",X"F4",X"F0",X"00",X"00",X"00",X"FF",X"98",X"88",X"8F",X"00",X"00",X"00",X"00",X"0F",
		X"88",X"89",X"99",X"8F",X"00",X"00",X"00",X"00",X"0F",X"FF",X"AA",X"77",X"F0",X"00",X"00",X"00",
		X"00",X"FE",X"BE",X"AA",X"77",X"F0",X"00",X"00",X"00",X"00",X"0F",X"F5",X"77",X"4F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F4",X"F7",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"75",
		X"4F",X"F0",X"00",X"00",X"00",X"00",X"F0",X"0F",X"55",X"55",X"EF",X"00",X"00",X"0F",X"FF",X"CF",
		X"FF",X"55",X"FF",X"5F",X"00",X"00",X"FC",X"CC",X"C5",X"EA",X"E5",X"EF",X"F5",X"F0",X"00",X"F9",
		X"99",X"5C",X"9E",X"45",X"EF",X"E5",X"F0",X"00",X"0F",X"FF",X"4E",X"95",X"4A",X"54",X"EF",X"05",
		X"00",X"00",X"0F",X"EC",X"9E",X"5A",X"EE",X"AE",X"E0",X"50",X"00",X"00",X"FF",X"FF",X"EB",X"FF",
		X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",X"FF",X"BF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"5B",X"EF",X"00",X"00",X"00",X"00",X"00",X"0F",X"4B",X"5F",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"98",X"88",X"8F",X"00",X"00",X"00",X"00",X"0F",X"88",X"89",X"99",X"8F",X"00",X"00",
		X"00",X"00",X"0F",X"FF",X"AA",X"77",X"F0",X"00",X"00",X"00",X"00",X"FE",X"BE",X"AA",X"77",X"F0",
		X"00",X"00",X"00",X"00",X"0F",X"F5",X"77",X"4F",X"FF",X"00",X"00",X"00",X"00",X"00",X"F4",X"F7",
		X"FF",X"5E",X"FF",X"00",X"00",X"00",X"00",X"0F",X"0F",X"77",X"54",X"5E",X"F0",X"00",X"00",X"FF",
		X"FC",X"FF",X"F5",X"5F",X"F5",X"EF",X"00",X"00",X"CC",X"CC",X"5E",X"AE",X"5E",X"FF",X"5F",X"00",
		X"00",X"99",X"95",X"C9",X"E4",X"5A",X"45",X"E0",X"E0",X"00",X"FF",X"F4",X"E9",X"55",X"5E",X"5E",
		X"FE",X"50",X"00",X"00",X"FE",X"C9",X"E5",X"EE",X"FF",X"00",X"E0",X"00",X"00",X"0F",X"FF",X"FE",
		X"B4",X"F0",X"EE",X"00",X"00",X"00",X"00",X"00",X"FB",X"FE",X"EF",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"BF",X"0F",X"F5",X"FF",X"00",X"00",X"00",X"00",X"FF",X"4B",X"F0",X"FF",X"55",X"F0",X"00",
		X"00",X"0F",X"BB",X"5F",X"0F",X"55",X"EF",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F8",X"88",X"F0",X"00",X"00",X"00",X"00",X"00",X"0F",X"88",X"88",
		X"8F",X"00",X"00",X"00",X"00",X"00",X"00",X"F9",X"99",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"B5",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"B7",X"4F",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"FF",X"7F",X"FF",X"00",X"00",X"00",X"00",X"00",X"FE",X"4E",X"7E",X"4E",X"F0",X"00",
		X"00",X"00",X"0F",X"E5",X"F5",X"E5",X"F5",X"EF",X"00",X"00",X"00",X"0F",X"5F",X"F5",X"55",X"FF",
		X"5F",X"00",X"00",X"00",X"0F",X"58",X"C8",X"55",X"E5",X"4F",X"00",X"00",X"00",X"00",X"F9",X"89",
		X"45",X"EE",X"5F",X"00",X"00",X"00",X"00",X"0F",X"EE",X"E4",X"5F",X"F0",X"00",X"00",X"00",X"00",
		X"0F",X"E5",X"55",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"4F",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"BF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"BF",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"B4",X"04",X"BF",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"88",X"89",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"99",X"98",X"88",X"F0",X"00",X"00",X"00",X"00",X"0F",X"77",X"AA",X"FF",X"F0",X"00",X"00",
		X"00",X"00",X"0F",X"77",X"AA",X"EB",X"EF",X"00",X"00",X"00",X"00",X"FF",X"F4",X"77",X"5F",X"F0",
		X"00",X"00",X"00",X"0F",X"E5",X"FF",X"7F",X"4F",X"00",X"00",X"00",X"00",X"F5",X"45",X"77",X"F0",
		X"F0",X"00",X"00",X"00",X"0F",X"5E",X"F5",X"5F",X"CF",X"FF",X"00",X"00",X"00",X"0F",X"5F",X"E5",
		X"E5",X"CC",X"CC",X"F0",X"00",X"00",X"0F",X"E5",X"EE",X"4E",X"59",X"99",X"F0",X"00",X"00",X"00",
		X"FE",X"45",X"E5",X"4F",X"FF",X"00",X"00",X"00",X"5E",X"EA",X"E5",X"AE",X"EF",X"00",X"00",X"00",
		X"05",X"0E",X"0F",X"F4",X"E5",X"F0",X"00",X"00",X"00",X"00",X"00",X"FF",X"BF",X"FF",X"5F",X"00",
		X"00",X"00",X"00",X"FF",X"B4",X"F0",X"00",X"F4",X"F0",X"00",X"00",X"0F",X"5B",X"FF",X"00",X"00",
		X"4E",X"4F",X"00",X"00",X"0F",X"4F",X"00",X"00",X"00",X"FF",X"FB",X"00",X"00",X"00",X"00",X"0F",
		X"88",X"88",X"9F",X"F0",X"00",X"00",X"00",X"00",X"0F",X"89",X"99",X"88",X"8F",X"00",X"00",X"00",
		X"00",X"00",X"F7",X"7A",X"AF",X"FF",X"00",X"00",X"00",X"00",X"00",X"F7",X"7A",X"AE",X"BE",X"F0",
		X"00",X"00",X"00",X"00",X"0F",X"47",X"75",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"F7",X"F4",
		X"F0",X"00",X"00",X"00",X"00",X"FF",X"45",X"7F",X"0F",X"00",X"00",X"00",X"00",X"0F",X"E5",X"55",
		X"5F",X"00",X"F0",X"00",X"00",X"00",X"0F",X"5F",X"F5",X"5F",X"FF",X"CF",X"FF",X"00",X"00",X"F5",
		X"FF",X"E5",X"EA",X"E5",X"CC",X"CC",X"F0",X"00",X"F5",X"EF",X"E5",X"4E",X"9C",X"59",X"99",X"F0",
		X"05",X"0F",X"E4",X"5A",X"45",X"9E",X"4F",X"FF",X"00",X"50",X"EE",X"AE",X"EA",X"5E",X"9C",X"EF",
		X"00",X"00",X"00",X"E0",X"FF",X"FB",X"EF",X"FF",X"F0",X"00",X"00",X"00",X"00",X"FF",X"BF",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"EB",X"5F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"5B",X"4F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"88",X"89",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"F8",X"99",X"98",X"88",X"F0",X"00",X"00",X"00",X"00",X"0F",X"77",X"AA",
		X"FF",X"F0",X"00",X"00",X"00",X"00",X"0F",X"77",X"AA",X"EB",X"EF",X"00",X"00",X"00",X"00",X"FF",
		X"F4",X"77",X"5F",X"F0",X"00",X"00",X"00",X"FF",X"E5",X"FF",X"7F",X"4F",X"00",X"00",X"00",X"0F",
		X"E5",X"45",X"77",X"F0",X"F0",X"00",X"00",X"00",X"FE",X"5F",X"F5",X"5F",X"FF",X"CF",X"FF",X"00",
		X"00",X"F5",X"FF",X"E5",X"EA",X"E5",X"CC",X"CC",X"00",X"0E",X"0E",X"54",X"A5",X"4E",X"9C",X"59",
		X"99",X"00",X"05",X"EF",X"E5",X"E5",X"55",X"9E",X"4F",X"FF",X"00",X"0E",X"00",X"FF",X"EE",X"5E",
		X"9C",X"EF",X"00",X"00",X"00",X"EE",X"0F",X"4B",X"EF",X"FF",X"F0",X"00",X"00",X"00",X"00",X"FE",
		X"EF",X"BF",X"00",X"00",X"00",X"00",X"00",X"FF",X"5F",X"F0",X"FB",X"F0",X"00",X"00",X"00",X"0F",
		X"55",X"FF",X"0F",X"B4",X"FF",X"00",X"00",X"00",X"00",X"FE",X"55",X"F0",X"F5",X"BB",X"F0",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"28",X"43",X"29",X"20",X"31",X"39",
		X"38",X"34",X"2C",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",
		X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
