library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity turkey_shoot_bank_b is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of turkey_shoot_bank_b is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"28",X"43",X"29",X"20",X"31",X"39",
		X"38",X"34",X"2C",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",
		X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"BD",X"F0",X"C4",
		X"BD",X"47",X"03",X"BD",X"40",X"2D",X"0F",X"6C",X"39",X"34",X"02",X"86",X"04",X"20",X"04",X"34",
		X"02",X"86",X"08",X"BA",X"C9",X"88",X"20",X"0D",X"34",X"02",X"86",X"FB",X"20",X"04",X"34",X"02",
		X"86",X"F7",X"B4",X"C9",X"88",X"B7",X"C9",X"88",X"35",X"82",X"0F",X"9B",X"96",X"50",X"84",X"C3",
		X"85",X"02",X"27",X"02",X"8A",X"10",X"D6",X"4E",X"C5",X"80",X"27",X"04",X"8A",X"24",X"03",X"9B",
		X"0D",X"E7",X"27",X"04",X"84",X"F0",X"9A",X"E8",X"1F",X"89",X"53",X"94",X"6C",X"D7",X"6C",X"97",
		X"41",X"39",X"34",X"07",X"1A",X"50",X"96",X"63",X"26",X"16",X"CC",X"06",X"05",X"97",X"63",X"D7",
		X"B3",X"96",X"50",X"D6",X"9D",X"27",X"02",X"8A",X"10",X"84",X"F7",X"B7",X"C9",X"86",X"97",X"50",
		X"35",X"87",X"86",X"02",X"34",X"01",X"1A",X"50",X"97",X"B3",X"96",X"50",X"84",X"F7",X"B7",X"C9",
		X"86",X"97",X"50",X"35",X"81",X"34",X"01",X"1A",X"50",X"96",X"64",X"26",X"0D",X"86",X"4B",X"97",
		X"64",X"96",X"50",X"8A",X"20",X"B7",X"C9",X"86",X"97",X"50",X"35",X"81",X"96",X"50",X"84",X"FB",
		X"B7",X"C9",X"86",X"0F",X"42",X"39",X"96",X"50",X"8A",X"04",X"B7",X"C9",X"86",X"39",X"D6",X"63",
		X"27",X"0B",X"0A",X"63",X"26",X"07",X"96",X"50",X"84",X"EF",X"B7",X"C9",X"86",X"D6",X"B3",X"27",
		X"0B",X"0A",X"B3",X"26",X"07",X"96",X"50",X"8A",X"08",X"B7",X"C9",X"86",X"D6",X"64",X"27",X"0B",
		X"0A",X"64",X"26",X"07",X"96",X"50",X"84",X"DF",X"B7",X"C9",X"86",X"39",X"96",X"39",X"27",X"02",
		X"0A",X"39",X"96",X"42",X"27",X"12",X"0A",X"42",X"26",X"0E",X"BD",X"00",X"CC",X"8E",X"70",X"75",
		X"BD",X"6F",X"D3",X"8E",X"EC",X"D5",X"9F",X"1D",X"39",X"96",X"41",X"85",X"40",X"26",X"05",X"85",
		X"80",X"26",X"08",X"39",X"C6",X"01",X"8E",X"A9",X"30",X"20",X"05",X"C6",X"02",X"8E",X"A9",X"33",
		X"D7",X"2C",X"96",X"8C",X"26",X"0A",X"B6",X"A9",X"43",X"90",X"2C",X"25",X"E6",X"B7",X"A9",X"43",
		X"86",X"01",X"BD",X"7E",X"EA",X"8E",X"A9",X"36",X"96",X"2C",X"BD",X"7E",X"EA",X"B6",X"A9",X"02",
		X"D6",X"2C",X"3D",X"1F",X"98",X"8E",X"A9",X"2D",X"BD",X"7E",X"EA",X"BD",X"DA",X"7F",X"0A",X"2C",
		X"0F",X"6C",X"7F",X"AA",X"60",X"7E",X"D4",X"02",X"39",X"1A",X"50",X"BD",X"E0",X"EC",X"C6",X"0C",
		X"BD",X"E5",X"61",X"1C",X"AF",X"8E",X"04",X"E0",X"BD",X"F5",X"42",X"8E",X"04",X"E6",X"BD",X"F5",
		X"4F",X"8E",X"04",X"EC",X"BD",X"F5",X"4F",X"8E",X"04",X"F2",X"BD",X"F5",X"4F",X"8E",X"00",X"17",
		X"BF",X"A5",X"C2",X"8E",X"00",X"A9",X"BF",X"A5",X"C8",X"CC",X"00",X"00",X"FD",X"A5",X"D5",X"FD",
		X"A5",X"D7",X"FD",X"A5",X"D9",X"FD",X"A5",X"DB",X"FD",X"A5",X"DD",X"FD",X"A5",X"DF",X"86",X"0F",
		X"B7",X"A5",X"D4",X"C6",X"33",X"BD",X"02",X"D7",X"7A",X"A5",X"D4",X"2C",X"F6",X"7F",X"A5",X"D4",
		X"C6",X"11",X"BD",X"D0",X"2D",X"86",X"04",X"BD",X"E0",X"76",X"BD",X"03",X"20",X"86",X"14",X"B7",
		X"A5",X"E3",X"86",X"FF",X"C6",X"40",X"D5",X"41",X"26",X"36",X"C6",X"01",X"D5",X"41",X"26",X"6C",
		X"40",X"C6",X"80",X"D5",X"41",X"26",X"29",X"C6",X"02",X"D5",X"41",X"26",X"5F",X"BD",X"E5",X"1F",
		X"96",X"60",X"27",X"DE",X"7E",X"03",X"3D",X"BD",X"E5",X"1F",X"96",X"50",X"B4",X"A5",X"E2",X"26",
		X"04",X"32",X"62",X"20",X"C8",X"7A",X"A5",X"E3",X"2C",X"ED",X"86",X"0A",X"B7",X"A5",X"E3",X"39",
		X"F7",X"A5",X"E2",X"B7",X"A5",X"E1",X"BB",X"A5",X"D4",X"2B",X"2A",X"81",X"0F",X"22",X"26",X"F6",
		X"A9",X"06",X"27",X"0E",X"81",X"04",X"26",X"04",X"8B",X"06",X"20",X"06",X"81",X"09",X"26",X"02",
		X"80",X"06",X"B7",X"A5",X"D4",X"BD",X"02",X"C9",X"C6",X"33",X"BD",X"D0",X"2D",X"BD",X"03",X"20",
		X"C6",X"11",X"BD",X"D0",X"2D",X"8D",X"B0",X"B6",X"A5",X"E1",X"20",X"CA",X"F7",X"A5",X"E2",X"B7",
		X"A5",X"E1",X"EC",X"D8",X"06",X"FB",X"A5",X"E1",X"2B",X"48",X"E1",X"48",X"24",X"44",X"1F",X"98",
		X"AE",X"44",X"27",X"02",X"A6",X"85",X"ED",X"D8",X"06",X"86",X"11",X"8D",X"3D",X"B6",X"A5",X"D4",
		X"81",X"03",X"26",X"28",X"B6",X"A9",X"06",X"27",X"23",X"4A",X"C6",X"07",X"3D",X"8E",X"04",X"89",
		X"3A",X"7C",X"A5",X"D4",X"BD",X"03",X"20",X"A6",X"80",X"2B",X"09",X"A7",X"D8",X"06",X"86",X"33",
		X"8D",X"18",X"20",X"ED",X"86",X"03",X"B7",X"A5",X"D4",X"BD",X"03",X"20",X"BD",X"DA",X"65",X"BD",
		X"DB",X"41",X"BD",X"02",X"07",X"B6",X"A5",X"E1",X"20",X"A8",X"34",X"10",X"8D",X"0B",X"C6",X"00",
		X"BD",X"D0",X"33",X"1F",X"89",X"8D",X"20",X"35",X"90",X"34",X"02",X"B6",X"A5",X"C4",X"8B",X"0C",
		X"B1",X"CB",X"E0",X"22",X"FB",X"35",X"82",X"F7",X"A5",X"C5",X"8D",X"44",X"AE",X"40",X"BF",X"A5",
		X"C0",X"8E",X"A5",X"C0",X"BD",X"F5",X"4F",X"F7",X"A5",X"CB",X"AE",X"42",X"27",X"08",X"EC",X"D8",
		X"06",X"58",X"AE",X"85",X"26",X"20",X"E6",X"D8",X"06",X"4F",X"BD",X"65",X"F9",X"8E",X"A5",X"CC",
		X"1F",X"98",X"BD",X"4B",X"4E",X"A6",X"1F",X"81",X"20",X"26",X"04",X"86",X"30",X"A7",X"1F",X"86",
		X"FF",X"A7",X"84",X"8E",X"A5",X"CC",X"BF",X"A5",X"C6",X"8E",X"A5",X"C6",X"BD",X"F5",X"4F",X"39",
		X"34",X"06",X"CE",X"03",X"93",X"B6",X"A5",X"D4",X"C6",X"09",X"3D",X"33",X"CB",X"B6",X"A5",X"D4",
		X"C6",X"0A",X"3D",X"CB",X"29",X"F7",X"A5",X"C4",X"F7",X"A5",X"CA",X"35",X"86",X"0F",X"60",X"7F",
		X"A5",X"E4",X"BD",X"E0",X"EC",X"86",X"04",X"BD",X"E0",X"76",X"B6",X"A5",X"D5",X"27",X"08",X"BD",
		X"DA",X"CC",X"8E",X"09",X"E1",X"8D",X"35",X"B6",X"A5",X"D7",X"27",X"08",X"BD",X"DA",X"DF",X"8E",
		X"09",X"DB",X"8D",X"28",X"B6",X"A5",X"D9",X"27",X"08",X"BD",X"DA",X"F8",X"8E",X"09",X"D5",X"8D",
		X"1B",X"B6",X"A5",X"E4",X"27",X"0D",X"86",X"F0",X"34",X"02",X"BD",X"E5",X"1F",X"6A",X"E4",X"26",
		X"F9",X"35",X"02",X"B6",X"A5",X"DB",X"27",X"03",X"BD",X"F2",X"C9",X"39",X"7C",X"A5",X"E4",X"BD",
		X"F5",X"42",X"39",X"05",X"94",X"04",X"25",X"04",X"4D",X"A9",X"00",X"14",X"05",X"A5",X"04",X"61",
		X"04",X"69",X"A9",X"02",X"04",X"05",X"C0",X"04",X"6D",X"00",X"00",X"A9",X"04",X"02",X"05",X"DF",
		X"04",X"75",X"00",X"00",X"A9",X"06",X"0A",X"05",X"F1",X"00",X"00",X"00",X"00",X"A9",X"08",X"63",
		X"06",X"03",X"00",X"00",X"00",X"00",X"A9",X"0A",X"63",X"06",X"17",X"00",X"00",X"00",X"00",X"A9",
		X"0C",X"63",X"06",X"2A",X"00",X"00",X"00",X"00",X"A9",X"0E",X"63",X"06",X"46",X"00",X"00",X"00",
		X"00",X"A9",X"10",X"63",X"06",X"68",X"00",X"00",X"00",X"00",X"A9",X"12",X"63",X"06",X"87",X"04",
		X"C8",X"00",X"00",X"A9",X"14",X"0A",X"05",X"D4",X"04",X"71",X"00",X"00",X"A9",X"18",X"02",X"06",
		X"9A",X"04",X"DC",X"00",X"00",X"A5",X"D5",X"02",X"06",X"B3",X"04",X"DC",X"00",X"00",X"A5",X"D7",
		X"02",X"06",X"CC",X"04",X"DC",X"00",X"00",X"A5",X"D9",X"02",X"06",X"E3",X"04",X"DC",X"00",X"00",
		X"A5",X"DB",X"02",X"00",X"00",X"06",X"EE",X"07",X"06",X"07",X"0C",X"07",X"12",X"07",X"18",X"07",
		X"1E",X"07",X"24",X"07",X"38",X"07",X"3E",X"07",X"4C",X"07",X"52",X"07",X"64",X"07",X"6A",X"07",
		X"7D",X"07",X"83",X"07",X"9C",X"07",X"A2",X"07",X"A8",X"07",X"AE",X"07",X"B4",X"00",X"05",X"0A",
		X"0F",X"14",X"19",X"1E",X"23",X"28",X"2D",X"32",X"37",X"3C",X"41",X"46",X"4B",X"50",X"55",X"5A",
		X"5F",X"07",X"C5",X"07",X"DF",X"07",X"F1",X"00",X"00",X"02",X"03",X"04",X"05",X"09",X"B7",X"09",
		X"B3",X"09",X"B7",X"09",X"B3",X"08",X"0A",X"08",X"28",X"08",X"40",X"08",X"55",X"08",X"6F",X"08",
		X"82",X"08",X"9A",X"08",X"AC",X"08",X"C0",X"08",X"CD",X"01",X"04",X"01",X"02",X"04",X"00",X"FF",
		X"06",X"00",X"01",X"01",X"00",X"00",X"FF",X"01",X"04",X"01",X"01",X"00",X"00",X"FF",X"01",X"10",
		X"06",X"02",X"00",X"00",X"FF",X"01",X"04",X"01",X"02",X"00",X"00",X"FF",X"01",X"00",X"04",X"01",
		X"00",X"00",X"FF",X"01",X"00",X"02",X"01",X"00",X"00",X"FF",X"01",X"00",X"02",X"02",X"00",X"00",
		X"FF",X"01",X"04",X"01",X"01",X"00",X"00",X"FF",X"08",X"DD",X"08",X"F5",X"09",X"09",X"09",X"1C",
		X"09",X"2A",X"09",X"41",X"09",X"53",X"09",X"6F",X"09",X"82",X"09",X"9A",X"09",X"B7",X"09",X"BB",
		X"04",X"F8",X"00",X"62",X"16",X"11",X"05",X"1F",X"00",X"1C",X"CE",X"11",X"05",X"5B",X"00",X"22",
		X"D6",X"11",X"05",X"09",X"00",X"68",X"E4",X"22",X"47",X"41",X"4D",X"45",X"20",X"41",X"44",X"4A",
		X"55",X"53",X"54",X"4D",X"45",X"4E",X"54",X"53",X"FF",X"50",X"52",X"45",X"53",X"53",X"20",X"41",
		X"44",X"56",X"41",X"4E",X"43",X"45",X"20",X"54",X"4F",X"20",X"45",X"58",X"49",X"54",X"FF",X"3C",
		X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"31",X"20",X"53",X"54",X"41",X"52",X"54",X"3E",X"20",
		X"54",X"4F",X"20",X"4D",X"4F",X"56",X"45",X"20",X"55",X"50",X"20",X"2D",X"20",X"3C",X"50",X"4C",
		X"41",X"59",X"45",X"52",X"20",X"32",X"20",X"53",X"54",X"41",X"52",X"54",X"3E",X"20",X"54",X"4F",
		X"20",X"4D",X"4F",X"56",X"45",X"20",X"44",X"4F",X"57",X"4E",X"FF",X"3C",X"47",X"4F",X"42",X"42",
		X"4C",X"45",X"3E",X"20",X"54",X"4F",X"20",X"49",X"4E",X"43",X"52",X"45",X"41",X"53",X"45",X"20",
		X"56",X"41",X"4C",X"55",X"45",X"20",X"2D",X"20",X"3C",X"47",X"52",X"45",X"4E",X"41",X"44",X"45",
		X"3E",X"20",X"54",X"4F",X"20",X"44",X"45",X"43",X"52",X"45",X"41",X"53",X"45",X"20",X"56",X"41",
		X"4C",X"55",X"45",X"FF",X"45",X"58",X"54",X"52",X"41",X"20",X"46",X"4F",X"57",X"4C",X"20",X"45",
		X"56",X"45",X"52",X"59",X"FF",X"4D",X"49",X"53",X"53",X"49",X"4F",X"4E",X"53",X"20",X"46",X"4F",
		X"52",X"20",X"31",X"20",X"43",X"52",X"45",X"44",X"49",X"54",X"20",X"47",X"41",X"4D",X"45",X"FF",
		X"41",X"54",X"54",X"52",X"41",X"43",X"54",X"20",X"4D",X"4F",X"44",X"45",X"20",X"53",X"4F",X"55",
		X"4E",X"44",X"53",X"FF",X"47",X"55",X"4E",X"20",X"52",X"45",X"43",X"4F",X"49",X"4C",X"FF",X"50",
		X"52",X"49",X"43",X"49",X"4E",X"47",X"20",X"53",X"45",X"4C",X"45",X"43",X"54",X"49",X"4F",X"4E",
		X"FF",X"20",X"20",X"4C",X"45",X"46",X"54",X"20",X"53",X"4C",X"4F",X"54",X"20",X"55",X"4E",X"49",
		X"54",X"53",X"FF",X"20",X"20",X"43",X"45",X"4E",X"54",X"45",X"52",X"20",X"53",X"4C",X"4F",X"54",
		X"20",X"55",X"4E",X"49",X"54",X"53",X"FF",X"20",X"20",X"52",X"49",X"47",X"48",X"54",X"20",X"53",
		X"4C",X"4F",X"54",X"20",X"55",X"4E",X"49",X"54",X"53",X"FF",X"20",X"20",X"55",X"4E",X"49",X"54",
		X"53",X"20",X"52",X"45",X"51",X"55",X"49",X"52",X"45",X"44",X"20",X"46",X"4F",X"52",X"20",X"43",
		X"52",X"45",X"44",X"49",X"54",X"FF",X"20",X"20",X"55",X"4E",X"49",X"54",X"53",X"20",X"52",X"45",
		X"51",X"55",X"49",X"52",X"45",X"44",X"20",X"46",X"4F",X"52",X"20",X"42",X"4F",X"4E",X"55",X"53",
		X"20",X"43",X"52",X"45",X"44",X"49",X"54",X"FF",X"20",X"20",X"4D",X"49",X"4E",X"49",X"4D",X"55",
		X"4D",X"20",X"55",X"4E",X"49",X"54",X"53",X"20",X"46",X"4F",X"52",X"20",X"41",X"4E",X"59",X"20",
		X"43",X"52",X"45",X"44",X"49",X"54",X"FF",X"44",X"49",X"46",X"46",X"49",X"43",X"55",X"4C",X"54",
		X"59",X"20",X"4F",X"46",X"20",X"50",X"4C",X"41",X"59",X"FF",X"52",X"45",X"53",X"54",X"4F",X"52",
		X"45",X"20",X"46",X"41",X"43",X"54",X"4F",X"52",X"59",X"20",X"53",X"45",X"54",X"54",X"49",X"4E",
		X"47",X"53",X"FF",X"43",X"4C",X"45",X"41",X"52",X"20",X"42",X"4F",X"4F",X"4B",X"4B",X"45",X"45",
		X"50",X"49",X"4E",X"47",X"20",X"54",X"4F",X"54",X"41",X"4C",X"53",X"FF",X"48",X"49",X"47",X"48",
		X"20",X"53",X"43",X"4F",X"52",X"45",X"20",X"54",X"41",X"42",X"4C",X"45",X"20",X"52",X"45",X"53",
		X"45",X"54",X"FF",X"41",X"55",X"54",X"4F",X"20",X"43",X"59",X"43",X"4C",X"45",X"FF",X"20",X"30",
		X"20",X"20",X"20",X"20",X"4E",X"4F",X"20",X"45",X"58",X"54",X"52",X"41",X"20",X"4D",X"49",X"53",
		X"53",X"49",X"4F",X"4E",X"53",X"FF",X"20",X"35",X"30",X"30",X"30",X"FF",X"31",X"30",X"30",X"30",
		X"30",X"FF",X"31",X"35",X"30",X"30",X"30",X"FF",X"32",X"30",X"30",X"30",X"30",X"FF",X"32",X"35",
		X"30",X"30",X"30",X"FF",X"33",X"30",X"30",X"30",X"30",X"20",X"45",X"58",X"54",X"52",X"41",X"20",
		X"4C",X"49",X"42",X"45",X"52",X"41",X"4C",X"FF",X"33",X"35",X"30",X"30",X"30",X"FF",X"34",X"30",
		X"30",X"30",X"30",X"20",X"4C",X"49",X"42",X"45",X"52",X"41",X"4C",X"FF",X"34",X"35",X"30",X"30",
		X"30",X"FF",X"35",X"30",X"30",X"30",X"30",X"20",X"52",X"45",X"43",X"4F",X"4D",X"4D",X"45",X"4E",
		X"44",X"45",X"44",X"FF",X"35",X"35",X"30",X"30",X"30",X"FF",X"36",X"30",X"30",X"30",X"30",X"20",
		X"43",X"4F",X"4E",X"53",X"45",X"52",X"56",X"41",X"54",X"49",X"56",X"45",X"FF",X"36",X"35",X"30",
		X"30",X"30",X"FF",X"37",X"30",X"30",X"30",X"30",X"20",X"45",X"58",X"54",X"52",X"41",X"20",X"43",
		X"4F",X"4E",X"53",X"45",X"52",X"56",X"41",X"54",X"49",X"56",X"45",X"FF",X"37",X"35",X"30",X"30",
		X"30",X"FF",X"38",X"30",X"30",X"30",X"30",X"FF",X"38",X"35",X"30",X"30",X"30",X"FF",X"39",X"30",
		X"30",X"30",X"30",X"FF",X"39",X"35",X"30",X"30",X"30",X"FF",X"20",X"55",X"4E",X"4C",X"49",X"4D",
		X"49",X"54",X"45",X"44",X"FF",X"20",X"32",X"20",X"20",X"20",X"20",X"48",X"49",X"47",X"48",X"20",
		X"56",X"4F",X"4C",X"55",X"4D",X"45",X"20",X"41",X"52",X"43",X"41",X"44",X"45",X"53",X"FF",X"20",
		X"33",X"20",X"20",X"20",X"20",X"52",X"45",X"43",X"4F",X"4D",X"4D",X"45",X"4E",X"44",X"45",X"44",
		X"FF",X"20",X"34",X"20",X"20",X"20",X"20",X"46",X"4F",X"52",X"20",X"57",X"45",X"41",X"4B",X"45",
		X"52",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"FF",X"20",X"30",X"20",X"20",X"20",X"20",
		X"43",X"55",X"53",X"54",X"4F",X"4D",X"20",X"2D",X"20",X"28",X"41",X"44",X"4A",X"55",X"53",X"54",
		X"20",X"42",X"45",X"4C",X"4F",X"57",X"29",X"FF",X"20",X"31",X"20",X"20",X"20",X"20",X"31",X"2F",
		X"46",X"49",X"46",X"54",X"59",X"20",X"20",X"33",X"2F",X"44",X"4F",X"4C",X"4C",X"41",X"52",X"FF",
		X"20",X"32",X"20",X"20",X"20",X"20",X"31",X"2F",X"31",X"20",X"44",X"4D",X"20",X"20",X"36",X"2F",
		X"35",X"20",X"44",X"4D",X"FF",X"20",X"33",X"20",X"20",X"20",X"20",X"31",X"2F",X"51",X"55",X"41",
		X"52",X"54",X"45",X"52",X"20",X"20",X"34",X"2F",X"44",X"4F",X"4C",X"4C",X"41",X"52",X"FF",X"20",
		X"34",X"20",X"20",X"20",X"20",X"31",X"2F",X"32",X"20",X"46",X"20",X"20",X"33",X"2F",X"35",X"20",
		X"46",X"FF",X"20",X"35",X"20",X"20",X"20",X"20",X"31",X"2F",X"46",X"49",X"46",X"54",X"59",X"20",
		X"20",X"32",X"2F",X"44",X"4F",X"4C",X"4C",X"41",X"52",X"FF",X"20",X"36",X"20",X"20",X"20",X"20",
		X"31",X"2F",X"32",X"35",X"20",X"20",X"34",X"2F",X"31",X"20",X"47",X"FF",X"20",X"37",X"20",X"20",
		X"20",X"20",X"31",X"2F",X"35",X"20",X"46",X"20",X"20",X"32",X"2F",X"31",X"30",X"20",X"46",X"FF",
		X"20",X"38",X"20",X"20",X"20",X"20",X"31",X"2F",X"31",X"30",X"20",X"46",X"FF",X"20",X"39",X"20",
		X"20",X"20",X"20",X"46",X"52",X"45",X"45",X"20",X"50",X"4C",X"41",X"59",X"FF",X"20",X"30",X"20",
		X"20",X"20",X"20",X"45",X"58",X"54",X"52",X"45",X"4D",X"45",X"4C",X"59",X"20",X"4C",X"49",X"42",
		X"45",X"52",X"41",X"4C",X"FF",X"20",X"31",X"20",X"20",X"20",X"20",X"45",X"58",X"54",X"52",X"41",
		X"20",X"4C",X"49",X"42",X"45",X"52",X"41",X"4C",X"FF",X"20",X"32",X"20",X"20",X"20",X"20",X"56",
		X"45",X"52",X"59",X"20",X"4C",X"49",X"42",X"45",X"52",X"41",X"4C",X"FF",X"20",X"33",X"20",X"20",
		X"20",X"20",X"4C",X"49",X"42",X"45",X"52",X"41",X"4C",X"FF",X"20",X"34",X"20",X"20",X"20",X"20",
		X"53",X"4F",X"4D",X"45",X"57",X"48",X"41",X"54",X"20",X"4C",X"49",X"42",X"45",X"52",X"41",X"4C",
		X"FF",X"20",X"35",X"20",X"20",X"20",X"20",X"52",X"45",X"43",X"4F",X"4D",X"4D",X"45",X"4E",X"44",
		X"45",X"44",X"FF",X"20",X"36",X"20",X"20",X"20",X"20",X"53",X"4F",X"4D",X"45",X"57",X"48",X"41",
		X"54",X"20",X"43",X"4F",X"4E",X"53",X"45",X"52",X"56",X"41",X"54",X"49",X"56",X"45",X"FF",X"20",
		X"37",X"20",X"20",X"20",X"20",X"43",X"4F",X"4E",X"53",X"45",X"52",X"56",X"41",X"54",X"49",X"56",
		X"45",X"FF",X"20",X"38",X"20",X"20",X"20",X"20",X"56",X"45",X"52",X"59",X"20",X"43",X"4F",X"4E",
		X"53",X"45",X"52",X"56",X"41",X"54",X"49",X"56",X"45",X"FF",X"20",X"39",X"20",X"20",X"20",X"20",
		X"45",X"58",X"54",X"52",X"41",X"20",X"43",X"4F",X"4E",X"53",X"45",X"52",X"56",X"41",X"54",X"49",
		X"56",X"45",X"FF",X"59",X"45",X"53",X"FF",X"4E",X"4F",X"20",X"FF",X"59",X"45",X"53",X"20",X"20",
		X"20",X"41",X"44",X"56",X"41",X"4E",X"43",X"45",X"20",X"54",X"4F",X"20",X"41",X"43",X"54",X"49",
		X"56",X"41",X"54",X"45",X"FF",X"0A",X"1C",X"00",X"50",X"50",X"22",X"0A",X"01",X"00",X"44",X"64",
		X"33",X"09",X"E7",X"00",X"47",X"78",X"11",X"46",X"41",X"43",X"54",X"4F",X"52",X"59",X"20",X"53",
		X"45",X"54",X"54",X"49",X"4E",X"47",X"53",X"20",X"52",X"45",X"53",X"54",X"4F",X"52",X"45",X"44",
		X"FF",X"42",X"4F",X"4F",X"4B",X"4B",X"45",X"45",X"50",X"49",X"4E",X"47",X"20",X"54",X"4F",X"54",
		X"41",X"4C",X"53",X"20",X"43",X"4C",X"45",X"41",X"52",X"45",X"44",X"FF",X"48",X"49",X"47",X"48",
		X"20",X"53",X"43",X"4F",X"52",X"45",X"20",X"54",X"41",X"42",X"4C",X"45",X"20",X"52",X"45",X"53",
		X"45",X"54",X"FF",X"3B",X"F8",X"3A",X"B8",X"3A",X"C2",X"3A",X"CC",X"3A",X"D6",X"3A",X"E0",X"3A",
		X"EA",X"3A",X"F4",X"3A",X"FE",X"3B",X"08",X"3B",X"12",X"3B",X"1C",X"3B",X"26",X"3B",X"30",X"3B",
		X"3A",X"3B",X"44",X"3B",X"4E",X"3B",X"58",X"3B",X"62",X"3B",X"6C",X"3B",X"76",X"3B",X"80",X"3B",
		X"8A",X"3B",X"94",X"3B",X"9E",X"3B",X"A8",X"3B",X"B2",X"3B",X"BC",X"3B",X"C6",X"3B",X"D0",X"3B",
		X"DA",X"3B",X"E4",X"3B",X"EE",X"39",X"B4",X"39",X"BE",X"39",X"C8",X"39",X"D2",X"39",X"DC",X"39",
		X"E6",X"39",X"F0",X"39",X"FA",X"3A",X"04",X"3A",X"0E",X"3A",X"18",X"3A",X"22",X"3A",X"2C",X"3A",
		X"36",X"3A",X"40",X"3A",X"4A",X"3A",X"54",X"3A",X"5E",X"3A",X"68",X"3A",X"72",X"3A",X"7C",X"3A",
		X"86",X"3A",X"90",X"3A",X"9A",X"3A",X"A4",X"3A",X"AE",X"3C",X"02",X"3C",X"0C",X"3C",X"16",X"3C",
		X"20",X"3C",X"2A",X"34",X"01",X"1A",X"50",X"BD",X"E0",X"EC",X"BD",X"E1",X"10",X"86",X"FF",X"97",
		X"9C",X"86",X"01",X"BD",X"E0",X"76",X"C6",X"04",X"BD",X"E5",X"61",X"1C",X"AF",X"BD",X"E5",X"1F",
		X"8E",X"10",X"5A",X"BD",X"F5",X"CC",X"8E",X"D5",X"21",X"A6",X"84",X"BD",X"66",X"BC",X"AE",X"01",
		X"BD",X"33",X"1B",X"0F",X"9C",X"BD",X"E5",X"1F",X"8D",X"1B",X"26",X"76",X"B6",X"BC",X"2D",X"2A",
		X"F4",X"86",X"B4",X"B7",X"A5",X"E5",X"BD",X"E5",X"1F",X"8D",X"0A",X"26",X"65",X"7A",X"A5",X"E5",
		X"26",X"F4",X"7E",X"0B",X"AE",X"96",X"41",X"84",X"01",X"39",X"8D",X"0C",X"8D",X"13",X"BD",X"E5",
		X"1F",X"8E",X"10",X"9A",X"BD",X"F4",X"87",X"39",X"BD",X"E5",X"1F",X"7D",X"BC",X"2D",X"2A",X"F8",
		X"39",X"BD",X"E5",X"1F",X"83",X"00",X"01",X"26",X"F8",X"39",X"BD",X"F5",X"CC",X"8D",X"E9",X"39",
		X"8D",X"F8",X"86",X"2D",X"BD",X"0D",X"5E",X"39",X"BD",X"F4",X"22",X"86",X"1E",X"BD",X"0D",X"5E",
		X"30",X"07",X"BD",X"F5",X"42",X"86",X"5A",X"BD",X"0D",X"5E",X"CC",X"0E",X"02",X"BD",X"33",X"3E",
		X"BD",X"0D",X"81",X"86",X"01",X"BD",X"E0",X"76",X"39",X"BD",X"F5",X"CC",X"CC",X"00",X"F0",X"8D",
		X"A9",X"39",X"BD",X"33",X"46",X"86",X"FF",X"97",X"9C",X"BD",X"E0",X"EC",X"BD",X"0D",X"8B",X"8E",
		X"0D",X"A4",X"BD",X"F4",X"44",X"CC",X"10",X"00",X"CE",X"E3",X"4E",X"BD",X"33",X"23",X"8E",X"10",
		X"A0",X"8D",X"D6",X"8E",X"11",X"44",X"8D",X"D1",X"8E",X"11",X"EA",X"8D",X"CC",X"8E",X"12",X"7F",
		X"BD",X"0B",X"2A",X"86",X"3C",X"BD",X"0D",X"5E",X"8E",X"12",X"FC",X"8D",X"BC",X"CC",X"10",X"00",
		X"BD",X"33",X"3E",X"BD",X"E0",X"EC",X"0F",X"9C",X"BE",X"D5",X"22",X"BD",X"33",X"1B",X"BD",X"0D",
		X"77",X"86",X"01",X"BD",X"E0",X"76",X"8E",X"0D",X"CF",X"BD",X"0B",X"2A",X"BD",X"0D",X"65",X"8E",
		X"0E",X"39",X"BD",X"0B",X"30",X"CE",X"0E",X"9B",X"10",X"8E",X"A5",X"E6",X"8E",X"00",X"1C",X"BD",
		X"7F",X"33",X"4F",X"F6",X"A9",X"02",X"BD",X"65",X"F9",X"8E",X"A5",X"F6",X"BD",X"66",X"1A",X"8E",
		X"0E",X"95",X"BD",X"0B",X"2A",X"BD",X"0D",X"65",X"8E",X"0E",X"B7",X"BD",X"0B",X"2A",X"86",X"5A",
		X"BD",X"0D",X"5E",X"8E",X"10",X"45",X"86",X"01",X"BD",X"F4",X"22",X"86",X"3C",X"BD",X"0D",X"5E",
		X"8E",X"10",X"4C",X"86",X"05",X"BD",X"F4",X"22",X"86",X"3C",X"BD",X"0D",X"5E",X"8E",X"10",X"53",
		X"86",X"01",X"BD",X"F4",X"22",X"86",X"B4",X"BD",X"0D",X"5E",X"CC",X"0E",X"02",X"BD",X"33",X"3E",
		X"BD",X"0D",X"77",X"86",X"01",X"BD",X"E0",X"76",X"8E",X"0E",X"D3",X"BD",X"0B",X"2A",X"86",X"78",
		X"BD",X"0D",X"5E",X"8E",X"0E",X"F2",X"BD",X"0B",X"30",X"8E",X"0F",X"FE",X"86",X"01",X"BD",X"0B",
		X"38",X"8E",X"0F",X"08",X"BD",X"0B",X"30",X"8E",X"10",X"18",X"86",X"05",X"BD",X"0B",X"38",X"8E",
		X"0F",X"1F",X"BD",X"0B",X"30",X"8E",X"10",X"0B",X"86",X"01",X"BD",X"0B",X"38",X"8E",X"0F",X"35",
		X"BD",X"0B",X"30",X"8E",X"10",X"25",X"86",X"01",X"BD",X"0B",X"38",X"BD",X"0D",X"77",X"8E",X"0F",
		X"56",X"BD",X"0B",X"2A",X"0F",X"E8",X"86",X"FF",X"97",X"E7",X"CC",X"8F",X"CF",X"DD",X"E5",X"BD",
		X"43",X"5B",X"CE",X"0D",X"AB",X"BD",X"0D",X"58",X"BD",X"E5",X"1F",X"CC",X"FF",X"00",X"BD",X"0D",
		X"3F",X"81",X"60",X"22",X"F3",X"BD",X"0D",X"47",X"CC",X"FF",X"00",X"BD",X"0D",X"3F",X"81",X"40",
		X"22",X"F6",X"BD",X"0D",X"47",X"BD",X"0D",X"65",X"8E",X"0F",X"78",X"BD",X"0B",X"2A",X"CE",X"0D",
		X"B1",X"BD",X"0D",X"58",X"86",X"13",X"BD",X"0D",X"5E",X"CE",X"0D",X"B1",X"BD",X"0D",X"58",X"CC",
		X"01",X"00",X"BD",X"0D",X"3F",X"81",X"63",X"25",X"F6",X"BD",X"0D",X"4B",X"86",X"64",X"BD",X"0D",
		X"5E",X"BD",X"0D",X"65",X"8E",X"0F",X"99",X"BD",X"0B",X"2A",X"BD",X"0D",X"65",X"8E",X"0F",X"D0",
		X"BD",X"0B",X"2A",X"86",X"FF",X"97",X"96",X"CE",X"0D",X"BD",X"BD",X"0D",X"58",X"86",X"08",X"BD",
		X"0D",X"5E",X"CE",X"0D",X"B7",X"BD",X"0D",X"58",X"CC",X"00",X"00",X"DD",X"D9",X"CC",X"FF",X"00",
		X"BD",X"0D",X"3F",X"81",X"20",X"22",X"F6",X"86",X"80",X"BD",X"0D",X"5E",X"CC",X"01",X"00",X"BD",
		X"0D",X"3F",X"81",X"65",X"25",X"F6",X"BD",X"0D",X"47",X"86",X"1E",X"BD",X"0D",X"5E",X"FE",X"B0",
		X"19",X"FC",X"51",X"2B",X"ED",X"C8",X"14",X"6F",X"C8",X"1D",X"CC",X"00",X"B4",X"BD",X"0B",X"21",
		X"FE",X"B0",X"3D",X"BD",X"43",X"8C",X"0F",X"E7",X"0F",X"96",X"BD",X"33",X"46",X"35",X"81",X"BD",
		X"E5",X"1F",X"D3",X"E5",X"DD",X"E5",X"39",X"86",X"04",X"20",X"02",X"86",X"01",X"BD",X"E5",X"1F",
		X"97",X"E8",X"BD",X"E5",X"1F",X"0F",X"E8",X"39",X"37",X"36",X"BD",X"63",X"61",X"39",X"BD",X"E5",
		X"1F",X"4A",X"26",X"FA",X"39",X"86",X"3C",X"8D",X"F5",X"CC",X"03",X"0B",X"BD",X"33",X"3E",X"8D",
		X"06",X"86",X"01",X"BD",X"E0",X"76",X"39",X"BD",X"E5",X"1F",X"8E",X"0D",X"C3",X"BD",X"F4",X"87",
		X"39",X"BD",X"E5",X"1F",X"8E",X"0D",X"C9",X"BD",X"F4",X"87",X"39",X"8E",X"10",X"82",X"BD",X"F4",
		X"87",X"8E",X"10",X"88",X"BD",X"F4",X"87",X"8E",X"10",X"8E",X"BD",X"F4",X"87",X"8E",X"10",X"94",
		X"BD",X"F4",X"87",X"39",X"20",X"00",X"00",X"59",X"28",X"39",X"28",X"00",X"04",X"01",X"CC",X"8F",
		X"CC",X"00",X"04",X"8F",X"CC",X"01",X"CC",X"00",X"04",X"01",X"CC",X"60",X"CC",X"00",X"0C",X"8F",
		X"CC",X"60",X"CC",X"00",X"00",X"4D",X"54",X"47",X"60",X"00",X"00",X"4D",X"68",X"47",X"60",X"0D",
		X"D5",X"00",X"4F",X"54",X"DD",X"41",X"73",X"20",X"61",X"20",X"54",X"75",X"72",X"6B",X"65",X"79",
		X"20",X"54",X"65",X"72",X"6D",X"69",X"6E",X"61",X"74",X"6F",X"72",X"2C",X"5C",X"79",X"6F",X"75",
		X"20",X"77",X"69",X"6C",X"6C",X"20",X"62",X"65",X"20",X"67",X"69",X"76",X"65",X"6E",X"20",X"31",
		X"30",X"30",X"5C",X"6D",X"69",X"73",X"73",X"69",X"6F",X"6E",X"73",X"2E",X"20",X"20",X"41",X"6C",
		X"6C",X"20",X"74",X"75",X"72",X"6B",X"65",X"79",X"73",X"5C",X"6D",X"75",X"73",X"74",X"20",X"62",
		X"65",X"20",X"65",X"6C",X"69",X"6D",X"69",X"6E",X"61",X"74",X"65",X"64",X"20",X"74",X"6F",X"5C",
		X"73",X"75",X"63",X"63",X"65",X"65",X"64",X"2E",X"FF",X"0E",X"3F",X"00",X"52",X"54",X"DD",X"41",
		X"20",X"6D",X"69",X"73",X"73",X"69",X"6F",X"6E",X"20",X"69",X"73",X"20",X"22",X"66",X"6F",X"75",
		X"6C",X"65",X"64",X"5C",X"75",X"70",X"22",X"20",X"69",X"66",X"20",X"61",X"20",X"74",X"75",X"72",
		X"6B",X"65",X"79",X"20",X"65",X"73",X"2D",X"5C",X"63",X"61",X"70",X"65",X"73",X"2C",X"20",X"6F",
		X"72",X"20",X"61",X"6E",X"79",X"20",X"69",X"6E",X"6E",X"6F",X"63",X"65",X"6E",X"74",X"5C",X"62",
		X"79",X"73",X"74",X"61",X"6E",X"64",X"65",X"72",X"20",X"69",X"73",X"20",X"64",X"61",X"6D",X"61",
		X"67",X"65",X"64",X"2E",X"FF",X"A5",X"E6",X"00",X"67",X"90",X"BB",X"59",X"6F",X"75",X"20",X"61",
		X"72",X"65",X"20",X"61",X"6C",X"6C",X"6F",X"77",X"65",X"64",X"5C",X"33",X"20",X"66",X"6F",X"75",
		X"6C",X"20",X"75",X"70",X"73",X"2E",X"FF",X"0E",X"BD",X"00",X"55",X"54",X"DD",X"50",X"72",X"6F",
		X"74",X"65",X"63",X"74",X"20",X"74",X"68",X"65",X"73",X"65",X"20",X"70",X"65",X"6F",X"70",X"6C",
		X"65",X"3A",X"FF",X"0E",X"D9",X"00",X"4C",X"54",X"11",X"50",X"72",X"65",X"73",X"65",X"6E",X"74",
		X"69",X"6E",X"67",X"20",X"74",X"68",X"65",X"20",X"76",X"69",X"6C",X"6C",X"61",X"69",X"6E",X"73",
		X"3A",X"FF",X"0E",X"F8",X"00",X"67",X"6C",X"BB",X"54",X"68",X"65",X"20",X"74",X"68",X"75",X"67",
		X"20",X"74",X"75",X"72",X"6B",X"65",X"79",X"FF",X"0F",X"0E",X"00",X"64",X"6C",X"BB",X"54",X"68",
		X"65",X"20",X"70",X"69",X"6C",X"6F",X"74",X"20",X"74",X"75",X"72",X"6B",X"65",X"79",X"FF",X"0F",
		X"25",X"00",X"67",X"6C",X"BB",X"54",X"68",X"65",X"20",X"62",X"6F",X"73",X"73",X"20",X"74",X"75",
		X"72",X"6B",X"65",X"79",X"FF",X"0F",X"3B",X"00",X"6D",X"6C",X"BB",X"54",X"68",X"65",X"20",X"63",
		X"79",X"62",X"6F",X"72",X"67",X"20",X"2D",X"5C",X"6D",X"65",X"63",X"68",X"61",X"6E",X"6F",X"74",
		X"75",X"72",X"6B",X"65",X"79",X"FF",X"0F",X"5C",X"00",X"64",X"54",X"DD",X"53",X"69",X"67",X"68",
		X"74",X"20",X"79",X"6F",X"75",X"72",X"20",X"65",X"6E",X"65",X"6D",X"79",X"5C",X"61",X"6E",X"64",
		X"20",X"73",X"68",X"6F",X"6F",X"74",X"21",X"FF",X"0F",X"7E",X"00",X"64",X"54",X"DD",X"4C",X"61",
		X"75",X"6E",X"63",X"68",X"20",X"61",X"20",X"67",X"72",X"65",X"6E",X"61",X"64",X"65",X"5C",X"77",
		X"68",X"65",X"6E",X"20",X"6C",X"69",X"74",X"2E",X"FF",X"0F",X"9F",X"00",X"61",X"54",X"DD",X"47",
		X"4F",X"42",X"42",X"4C",X"45",X"20",X"62",X"75",X"74",X"74",X"6F",X"6E",X"20",X"6D",X"61",X"79",
		X"5C",X"62",X"65",X"20",X"75",X"73",X"65",X"64",X"20",X"6F",X"6E",X"6C",X"79",X"20",X"6F",X"6E",
		X"63",X"65",X"5C",X"70",X"65",X"72",X"20",X"6D",X"69",X"73",X"73",X"69",X"6F",X"6E",X"2E",X"FF",
		X"0F",X"D6",X"00",X"5B",X"54",X"DD",X"54",X"61",X"6B",X"65",X"20",X"63",X"61",X"72",X"65",X"66",
		X"75",X"6C",X"20",X"61",X"69",X"6D",X"20",X"69",X"66",X"5C",X"61",X"20",X"68",X"6F",X"73",X"74",
		X"61",X"67",X"65",X"20",X"69",X"73",X"20",X"74",X"61",X"6B",X"65",X"6E",X"2E",X"FF",X"63",X"05",
		X"00",X"88",X"95",X"0C",X"19",X"10",X"32",X"00",X"85",X"BA",X"DD",X"07",X"FC",X"00",X"89",X"93",
		X"0B",X"1B",X"10",X"38",X"00",X"85",X"BA",X"DD",X"20",X"2D",X"00",X"89",X"9D",X"0B",X"1A",X"10",
		X"32",X"00",X"85",X"BA",X"DD",X"46",X"45",X"00",X"89",X"90",X"0B",X"1E",X"10",X"3E",X"00",X"82",
		X"BA",X"DD",X"28",X"35",X"30",X"30",X"29",X"FF",X"28",X"37",X"35",X"30",X"29",X"FF",X"28",X"31",
		X"30",X"30",X"30",X"29",X"FF",X"25",X"0D",X"00",X"70",X"70",X"08",X"1A",X"2A",X"58",X"00",X"8E",
		X"71",X"07",X"19",X"2F",X"AA",X"00",X"AC",X"74",X"07",X"16",X"10",X"60",X"00",X"58",X"54",X"BB",
		X"5C",X"5C",X"50",X"72",X"65",X"73",X"73",X"20",X"47",X"52",X"45",X"4E",X"41",X"44",X"45",X"20",
		X"62",X"75",X"74",X"74",X"6F",X"6E",X"5C",X"66",X"6F",X"72",X"20",X"73",X"74",X"6F",X"72",X"79",
		X"2E",X"FF",X"E0",X"00",X"14",X"18",X"01",X"C8",X"0E",X"01",X"0F",X"18",X"01",X"C8",X"EE",X"00",
		X"14",X"18",X"7E",X"01",X"EE",X"00",X"14",X"E0",X"7E",X"01",X"00",X"00",X"28",X"64",X"69",X"6C",
		X"10",X"A6",X"00",X"32",X"64",X"88",X"54",X"68",X"65",X"20",X"79",X"65",X"61",X"72",X"20",X"69",
		X"73",X"20",X"31",X"39",X"38",X"39",X"2C",X"20",X"6F",X"6E",X"65",X"20",X"79",X"65",X"61",X"72",
		X"20",X"61",X"66",X"74",X"65",X"72",X"5C",X"74",X"68",X"65",X"20",X"67",X"72",X"65",X"61",X"74",
		X"20",X"67",X"6F",X"62",X"62",X"6C",X"65",X"20",X"62",X"6C",X"69",X"67",X"68",X"74",X"20",X"77",
		X"68",X"69",X"63",X"68",X"5C",X"70",X"6C",X"61",X"67",X"75",X"65",X"64",X"20",X"74",X"68",X"65",
		X"20",X"77",X"6F",X"72",X"6C",X"64",X"2E",X"20",X"20",X"4F",X"6E",X"65",X"20",X"74",X"68",X"69",
		X"72",X"64",X"20",X"6F",X"66",X"5C",X"65",X"61",X"72",X"74",X"68",X"27",X"73",X"20",X"70",X"6F",
		X"70",X"75",X"6C",X"61",X"63",X"65",X"20",X"77",X"61",X"73",X"20",X"74",X"72",X"61",X"6E",X"73",
		X"66",X"6F",X"72",X"6D",X"65",X"64",X"5C",X"69",X"6E",X"74",X"6F",X"20",X"74",X"75",X"72",X"6B",
		X"65",X"79",X"73",X"20",X"62",X"79",X"20",X"74",X"68",X"65",X"20",X"61",X"69",X"6C",X"6D",X"65",
		X"6E",X"74",X"2E",X"FF",X"11",X"4A",X"00",X"2C",X"64",X"88",X"54",X"68",X"65",X"20",X"73",X"69",
		X"64",X"65",X"20",X"65",X"66",X"66",X"65",X"63",X"74",X"20",X"6F",X"66",X"20",X"74",X"75",X"72",
		X"6B",X"65",X"79",X"20",X"74",X"72",X"61",X"6E",X"73",X"2D",X"5C",X"66",X"6F",X"72",X"6D",X"61",
		X"74",X"69",X"6F",X"6E",X"20",X"69",X"73",X"20",X"61",X"20",X"74",X"65",X"6E",X"64",X"65",X"6E",
		X"63",X"79",X"20",X"74",X"6F",X"77",X"61",X"72",X"64",X"5C",X"76",X"69",X"6F",X"6C",X"65",X"6E",
		X"63",X"65",X"20",X"61",X"6E",X"64",X"20",X"63",X"6F",X"6D",X"72",X"61",X"64",X"65",X"72",X"79",
		X"20",X"62",X"65",X"74",X"77",X"65",X"65",X"6E",X"5C",X"74",X"68",X"65",X"73",X"65",X"20",X"74",
		X"75",X"72",X"6B",X"65",X"79",X"73",X"20",X"74",X"6F",X"20",X"6F",X"72",X"67",X"61",X"6E",X"69",
		X"7A",X"65",X"20",X"66",X"6F",X"72",X"5C",X"72",X"61",X"62",X"62",X"6C",X"65",X"2D",X"72",X"6F",
		X"75",X"73",X"69",X"6E",X"67",X"20",X"69",X"6E",X"20",X"74",X"68",X"65",X"20",X"75",X"72",X"62",
		X"61",X"6E",X"20",X"61",X"72",X"65",X"61",X"73",X"2E",X"FF",X"11",X"F0",X"00",X"35",X"64",X"88",
		X"49",X"6E",X"20",X"46",X"65",X"62",X"72",X"75",X"61",X"72",X"79",X"20",X"6F",X"66",X"20",X"27",
		X"38",X"39",X"2C",X"20",X"61",X"20",X"67",X"72",X"6F",X"75",X"70",X"20",X"6F",X"66",X"5C",X"73",
		X"70",X"65",X"63",X"69",X"61",X"6C",X"6C",X"79",X"20",X"74",X"72",X"61",X"69",X"6E",X"65",X"64",
		X"20",X"61",X"67",X"65",X"6E",X"74",X"73",X"20",X"28",X"74",X"68",X"65",X"5C",X"54",X"75",X"72",
		X"6B",X"65",X"79",X"20",X"54",X"65",X"72",X"6D",X"69",X"6E",X"61",X"74",X"6F",X"72",X"73",X"29",
		X"20",X"77",X"61",X"73",X"20",X"66",X"6F",X"72",X"6D",X"65",X"64",X"5C",X"66",X"6F",X"72",X"20",
		X"74",X"68",X"65",X"20",X"73",X"6F",X"6C",X"65",X"20",X"74",X"61",X"73",X"6B",X"20",X"6F",X"66",
		X"20",X"64",X"65",X"73",X"74",X"72",X"6F",X"79",X"69",X"6E",X"67",X"5C",X"74",X"68",X"65",X"20",
		X"74",X"75",X"72",X"6B",X"65",X"79",X"20",X"6D",X"65",X"6E",X"61",X"63",X"65",X"2E",X"FF",X"12",
		X"85",X"00",X"38",X"64",X"88",X"41",X"73",X"20",X"61",X"20",X"74",X"65",X"72",X"6D",X"69",X"6E",
		X"61",X"74",X"6F",X"72",X"2C",X"20",X"79",X"6F",X"75",X"20",X"6D",X"75",X"73",X"74",X"20",X"62",
		X"65",X"5C",X"6D",X"65",X"6E",X"74",X"61",X"6C",X"6C",X"79",X"20",X"61",X"6E",X"64",X"20",X"70",
		X"68",X"79",X"73",X"69",X"63",X"61",X"6C",X"6C",X"79",X"20",X"70",X"72",X"65",X"2D",X"5C",X"70",
		X"61",X"72",X"65",X"64",X"20",X"66",X"6F",X"72",X"20",X"61",X"20",X"73",X"65",X"72",X"69",X"65",
		X"73",X"20",X"6F",X"66",X"20",X"6D",X"69",X"73",X"73",X"69",X"6F",X"6E",X"73",X"5C",X"63",X"6F",
		X"6D",X"70",X"6C",X"69",X"6D",X"65",X"6E",X"74",X"61",X"72",X"79",X"20",X"74",X"6F",X"20",X"79",
		X"6F",X"75",X"72",X"20",X"73",X"6B",X"69",X"6C",X"6C",X"73",X"2E",X"FF",X"13",X"02",X"00",X"38",
		X"A0",X"99",X"47",X"6F",X"6F",X"64",X"20",X"6C",X"75",X"63",X"6B",X"20",X"61",X"6E",X"64",X"20",
		X"73",X"74",X"72",X"65",X"6E",X"67",X"74",X"68",X"20",X"74",X"6F",X"20",X"79",X"6F",X"75",X"21",
		X"FF",X"39",X"34",X"76",X"CE",X"A6",X"90",X"EC",X"81",X"ED",X"44",X"A6",X"80",X"A7",X"43",X"EC",
		X"81",X"FD",X"A6",X"8D",X"EC",X"81",X"FD",X"A6",X"8A",X"48",X"A7",X"42",X"E7",X"41",X"A6",X"80",
		X"B7",X"A6",X"8F",X"10",X"AE",X"81",X"10",X"BF",X"A6",X"96",X"17",X"00",X"71",X"B6",X"A6",X"8E",
		X"A7",X"40",X"6F",X"41",X"8D",X"79",X"AF",X"44",X"B6",X"A6",X"8B",X"A7",X"41",X"A6",X"43",X"AB",
		X"41",X"A7",X"43",X"8D",X"49",X"8D",X"68",X"E7",X"43",X"B6",X"A6",X"8A",X"40",X"48",X"A7",X"42",
		X"AE",X"44",X"30",X"86",X"AF",X"44",X"6F",X"41",X"7A",X"A6",X"8E",X"B6",X"A6",X"8E",X"A7",X"40",
		X"8D",X"4D",X"AF",X"44",X"B6",X"A6",X"8B",X"40",X"A7",X"41",X"A6",X"43",X"AB",X"41",X"A7",X"43",
		X"8D",X"1C",X"8D",X"3B",X"E7",X"43",X"B6",X"A6",X"8A",X"48",X"A7",X"42",X"AE",X"44",X"30",X"86",
		X"AF",X"44",X"7A",X"A6",X"8E",X"8D",X"17",X"7A",X"A6",X"8F",X"26",X"A1",X"35",X"F6",X"6F",X"42",
		X"B6",X"A6",X"8D",X"4A",X"26",X"02",X"86",X"01",X"B7",X"A6",X"8D",X"A7",X"40",X"39",X"BE",X"A6",
		X"96",X"10",X"AE",X"81",X"26",X"05",X"AE",X"84",X"10",X"AE",X"81",X"BF",X"A6",X"96",X"39",X"EC",
		X"C4",X"34",X"06",X"EC",X"42",X"AE",X"44",X"20",X"04",X"30",X"86",X"EB",X"61",X"BF",X"A6",X"87",
		X"F7",X"A6",X"89",X"34",X"16",X"A6",X"A0",X"26",X"05",X"10",X"AE",X"A1",X"A6",X"A0",X"B7",X"A6",
		X"86",X"8E",X"A6",X"86",X"BD",X"F4",X"87",X"35",X"16",X"6A",X"E4",X"26",X"DC",X"32",X"61",X"35",
		X"82",X"CE",X"1A",X"C9",X"10",X"8E",X"A8",X"E2",X"8E",X"00",X"10",X"BD",X"7F",X"33",X"39",X"86",
		X"01",X"A7",X"C8",X"1F",X"6F",X"C8",X"57",X"BD",X"63",X"23",X"AF",X"C8",X"54",X"6F",X"C8",X"56",
		X"11",X"A3",X"88",X"54",X"26",X"0A",X"A6",X"88",X"56",X"2B",X"02",X"86",X"01",X"A7",X"C8",X"56",
		X"CC",X"1A",X"27",X"ED",X"C8",X"40",X"CC",X"00",X"00",X"A7",X"4E",X"A7",X"C8",X"1D",X"ED",X"C8",
		X"34",X"ED",X"C8",X"36",X"ED",X"C8",X"47",X"A7",X"C8",X"38",X"A7",X"C8",X"3A",X"A7",X"C8",X"42",
		X"A7",X"C8",X"44",X"A7",X"C8",X"45",X"A7",X"C8",X"4A",X"A7",X"C8",X"4B",X"ED",X"C8",X"4C",X"A7",
		X"C8",X"4E",X"A7",X"C8",X"50",X"A7",X"C8",X"51",X"A7",X"C8",X"52",X"A7",X"C8",X"53",X"A7",X"C8",
		X"58",X"A7",X"C8",X"59",X"A7",X"C8",X"4F",X"B6",X"A8",X"F2",X"A7",X"C8",X"3C",X"A7",X"C8",X"3B",
		X"8E",X"14",X"8F",X"AF",X"C8",X"3E",X"8E",X"14",X"8C",X"AF",X"4A",X"39",X"6E",X"D8",X"3E",X"A6",
		X"4E",X"27",X"28",X"AE",X"C8",X"4C",X"27",X"0C",X"CC",X"00",X"00",X"ED",X"88",X"4C",X"A7",X"88",
		X"4B",X"A7",X"88",X"4E",X"AE",X"C8",X"54",X"27",X"0E",X"A6",X"C8",X"56",X"27",X"09",X"CC",X"00",
		X"00",X"ED",X"88",X"54",X"A7",X"88",X"56",X"BD",X"30",X"7C",X"39",X"8E",X"16",X"64",X"AF",X"C8",
		X"3E",X"FC",X"A8",X"DA",X"6D",X"C8",X"4E",X"27",X"03",X"CC",X"02",X"00",X"FD",X"A8",X"DE",X"CC",
		X"00",X"00",X"B3",X"A8",X"DE",X"FD",X"A8",X"E0",X"EC",X"C8",X"14",X"ED",X"C8",X"5E",X"0D",X"39",
		X"27",X"1F",X"AE",X"C8",X"4C",X"27",X"12",X"CC",X"00",X"00",X"A7",X"C8",X"4E",X"ED",X"C8",X"4C",
		X"ED",X"88",X"4C",X"A7",X"88",X"4B",X"A7",X"88",X"4E",X"8E",X"00",X"00",X"AF",X"C8",X"36",X"20",
		X"7A",X"E0",X"C8",X"32",X"2A",X"01",X"50",X"C1",X"08",X"23",X"05",X"EC",X"C8",X"36",X"26",X"71",
		X"86",X"FF",X"A7",X"C8",X"53",X"6F",X"C8",X"58",X"EC",X"C8",X"14",X"E1",X"C8",X"32",X"25",X"3E",
		X"22",X"42",X"10",X"8E",X"00",X"00",X"A1",X"C8",X"30",X"25",X"49",X"22",X"42",X"A6",X"C8",X"1D",
		X"26",X"4C",X"86",X"FF",X"A7",X"C8",X"1D",X"BD",X"39",X"13",X"B6",X"A8",X"F2",X"A7",X"C8",X"3C",
		X"A6",X"C8",X"4B",X"27",X"14",X"AE",X"C8",X"4C",X"27",X"0F",X"A7",X"88",X"4B",X"A7",X"C8",X"4E",
		X"6F",X"C8",X"4B",X"8E",X"70",X"A9",X"BD",X"6F",X"D3",X"8E",X"00",X"00",X"20",X"19",X"10",X"BE",
		X"A8",X"E0",X"20",X"04",X"10",X"BE",X"A8",X"DE",X"A1",X"C8",X"30",X"25",X"07",X"27",X"EA",X"BE",
		X"A8",X"DE",X"20",X"03",X"BE",X"A8",X"E0",X"10",X"AF",X"C8",X"36",X"AF",X"C8",X"34",X"7E",X"1A",
		X"20",X"6F",X"C8",X"53",X"A6",X"C8",X"58",X"26",X"37",X"A6",X"C8",X"50",X"26",X"15",X"A6",X"C8",
		X"51",X"26",X"1A",X"A6",X"C8",X"14",X"A1",X"C8",X"30",X"22",X"04",X"8D",X"4E",X"20",X"49",X"8D",
		X"50",X"20",X"45",X"6A",X"C8",X"50",X"A6",X"C8",X"52",X"2D",X"0A",X"20",X"0D",X"6A",X"C8",X"51",
		X"A6",X"C8",X"52",X"2D",X"05",X"BE",X"A8",X"E0",X"20",X"03",X"BE",X"A8",X"DE",X"AF",X"C8",X"34",
		X"E6",X"C8",X"15",X"E1",X"C8",X"32",X"25",X"07",X"22",X"0A",X"8E",X"00",X"00",X"20",X"08",X"BE",
		X"A8",X"E0",X"20",X"03",X"BE",X"A8",X"DE",X"AF",X"C8",X"36",X"A6",X"C8",X"38",X"27",X"26",X"6F",
		X"C8",X"58",X"B6",X"A8",X"F2",X"A7",X"C8",X"3C",X"7E",X"1A",X"20",X"34",X"06",X"86",X"FF",X"20",
		X"03",X"34",X"06",X"4F",X"A7",X"C8",X"52",X"DC",X"D5",X"84",X"03",X"C4",X"03",X"C3",X"0A",X"02",
		X"ED",X"C8",X"50",X"35",X"86",X"A6",X"C8",X"58",X"26",X"1B",X"6C",X"C8",X"59",X"A6",X"C8",X"59",
		X"81",X"04",X"25",X"4D",X"6F",X"C8",X"59",X"6C",X"C8",X"58",X"6F",X"C8",X"3C",X"8E",X"70",X"AD",
		X"BD",X"6F",X"D3",X"20",X"3C",X"EC",X"C8",X"34",X"2B",X"07",X"27",X"0B",X"CC",X"00",X"40",X"20",
		X"03",X"CC",X"FF",X"C0",X"ED",X"C8",X"34",X"8E",X"1B",X"29",X"E6",X"C8",X"4E",X"27",X"03",X"8E",
		X"1B",X"3D",X"A6",X"C8",X"58",X"48",X"EC",X"86",X"E3",X"C8",X"36",X"ED",X"C8",X"36",X"6C",X"C8",
		X"58",X"A6",X"C8",X"58",X"81",X"0A",X"26",X"09",X"6F",X"C8",X"58",X"B6",X"A8",X"F2",X"A7",X"C8",
		X"3C",X"7E",X"1A",X"20",X"8E",X"18",X"A2",X"AF",X"C8",X"3E",X"A6",X"C8",X"30",X"E6",X"C8",X"32",
		X"BD",X"67",X"5E",X"A7",X"C8",X"38",X"27",X"08",X"A7",X"C8",X"16",X"8E",X"16",X"83",X"AF",X"4A",
		X"7E",X"1A",X"20",X"A6",X"C8",X"16",X"8E",X"1A",X"61",X"AE",X"86",X"A6",X"C8",X"30",X"E6",X"C8",
		X"32",X"10",X"A3",X"C8",X"5E",X"26",X"09",X"6D",X"C8",X"56",X"2D",X"04",X"1A",X"04",X"6E",X"84",
		X"1C",X"FB",X"6E",X"84",X"10",X"26",X"01",X"13",X"CC",X"14",X"30",X"7E",X"17",X"04",X"10",X"26",
		X"01",X"11",X"CC",X"26",X"30",X"20",X"4D",X"10",X"26",X"01",X"10",X"CC",X"46",X"30",X"20",X"44",
		X"10",X"26",X"00",X"FF",X"CC",X"6B",X"30",X"20",X"3B",X"10",X"26",X"00",X"EE",X"CC",X"83",X"30",
		X"20",X"32",X"10",X"26",X"00",X"DD",X"C6",X"A1",X"8E",X"1A",X"D9",X"20",X"2E",X"10",X"26",X"00",
		X"D2",X"C6",X"A1",X"8E",X"1A",X"F1",X"20",X"23",X"10",X"26",X"00",X"DF",X"C6",X"31",X"8E",X"1B",
		X"09",X"20",X"18",X"10",X"26",X"00",X"D4",X"C6",X"31",X"8E",X"1B",X"19",X"20",X"0D",X"CC",X"14",
		X"8C",X"ED",X"4A",X"39",X"8E",X"A8",X"E2",X"A7",X"01",X"A7",X"09",X"E7",X"45",X"20",X"60",X"6A",
		X"C8",X"1C",X"26",X"70",X"8E",X"A8",X"EA",X"20",X"56",X"6A",X"C8",X"1C",X"26",X"66",X"8E",X"1A",
		X"E1",X"20",X"4C",X"6A",X"C8",X"1C",X"26",X"5C",X"8E",X"1A",X"E9",X"20",X"42",X"6A",X"C8",X"1C",
		X"26",X"52",X"8E",X"1A",X"F9",X"20",X"38",X"6A",X"C8",X"1C",X"26",X"48",X"8E",X"1B",X"01",X"20",
		X"2E",X"10",X"26",X"01",X"07",X"0D",X"E4",X"10",X"26",X"01",X"01",X"8E",X"1A",X"A9",X"20",X"1F",
		X"10",X"26",X"01",X"0E",X"8E",X"1A",X"B9",X"20",X"16",X"10",X"26",X"00",X"FA",X"0D",X"E4",X"10",
		X"26",X"00",X"F4",X"8E",X"1A",X"A1",X"20",X"07",X"10",X"26",X"01",X"01",X"8E",X"1A",X"B1",X"EC",
		X"81",X"A7",X"C8",X"1C",X"E7",X"44",X"EC",X"81",X"ED",X"42",X"6C",X"4F",X"EC",X"81",X"ED",X"46",
		X"EC",X"84",X"ED",X"4A",X"39",X"6A",X"C8",X"1C",X"26",X"FA",X"8E",X"1A",X"C1",X"20",X"E0",X"6A",
		X"C8",X"1C",X"26",X"F0",X"8E",X"1B",X"11",X"20",X"D6",X"6A",X"C8",X"1C",X"26",X"E6",X"8E",X"1B",
		X"21",X"20",X"CC",X"27",X"E5",X"20",X"0C",X"27",X"E1",X"20",X"10",X"C1",X"EC",X"25",X"5D",X"C6",
		X"EC",X"20",X"3F",X"C1",X"B1",X"22",X"55",X"C6",X"B1",X"20",X"27",X"C1",X"39",X"25",X"04",X"C6",
		X"39",X"20",X"2F",X"C1",X"37",X"22",X"45",X"C6",X"37",X"20",X"17",X"C1",X"38",X"22",X"3D",X"C6",
		X"38",X"20",X"0F",X"C1",X"97",X"22",X"35",X"C6",X"98",X"8E",X"00",X"00",X"AF",X"C8",X"34",X"BD",
		X"39",X"2F",X"E7",X"C8",X"32",X"EC",X"C8",X"36",X"2A",X"22",X"CC",X"00",X"00",X"ED",X"C8",X"36",
		X"20",X"1A",X"E7",X"C8",X"32",X"EC",X"C8",X"36",X"2F",X"12",X"20",X"EE",X"C1",X"68",X"25",X"0C",
		X"C6",X"68",X"20",X"EE",X"C1",X"48",X"25",X"04",X"C6",X"48",X"20",X"E6",X"CC",X"14",X"8C",X"ED",
		X"4A",X"39",X"A7",X"C8",X"30",X"EC",X"C8",X"34",X"2A",X"F2",X"CC",X"00",X"00",X"ED",X"C8",X"34",
		X"20",X"EA",X"A7",X"C8",X"30",X"EC",X"C8",X"34",X"2F",X"E2",X"20",X"EE",X"81",X"24",X"22",X"DC",
		X"86",X"24",X"20",X"DE",X"81",X"70",X"25",X"D4",X"86",X"70",X"20",X"E6",X"81",X"1C",X"22",X"CC",
		X"86",X"1C",X"20",X"CE",X"81",X"75",X"25",X"C4",X"86",X"75",X"20",X"D6",X"BD",X"15",X"F1",X"81",
		X"25",X"22",X"B9",X"86",X"25",X"20",X"BB",X"BD",X"15",X"EB",X"81",X"6E",X"25",X"AE",X"86",X"6E",
		X"20",X"C0",X"BD",X"15",X"F1",X"81",X"28",X"22",X"A3",X"86",X"28",X"20",X"A5",X"BD",X"15",X"EB",
		X"81",X"6C",X"25",X"98",X"86",X"6C",X"20",X"AA",X"C6",X"10",X"E7",X"C8",X"14",X"E6",X"C8",X"32",
		X"E7",X"C8",X"15",X"C6",X"FF",X"E7",X"C8",X"1E",X"86",X"01",X"20",X"86",X"C6",X"80",X"E7",X"C8",
		X"14",X"E6",X"C8",X"32",X"E7",X"C8",X"15",X"C6",X"FF",X"E7",X"C8",X"1E",X"20",X"84",X"BD",X"38",
		X"52",X"39",X"8E",X"19",X"3F",X"AF",X"C8",X"3E",X"A6",X"C8",X"4E",X"27",X"06",X"AE",X"C8",X"4C",
		X"A7",X"88",X"4E",X"A6",X"C8",X"48",X"BB",X"A8",X"F3",X"A7",X"C8",X"48",X"24",X"0B",X"6C",X"C8",
		X"47",X"6A",X"C8",X"3C",X"2A",X"03",X"6F",X"C8",X"3C",X"A6",X"C8",X"53",X"26",X"08",X"EC",X"C8",
		X"36",X"E3",X"C8",X"32",X"20",X"30",X"EC",X"C8",X"36",X"2D",X"20",X"26",X"14",X"EC",X"C8",X"34",
		X"26",X"27",X"6C",X"C8",X"4A",X"A6",X"C8",X"4A",X"81",X"08",X"25",X"20",X"BD",X"39",X"2F",X"20",
		X"18",X"E3",X"C8",X"32",X"A1",X"C8",X"5F",X"22",X"0A",X"20",X"0B",X"E3",X"C8",X"32",X"A1",X"C8",
		X"5F",X"24",X"03",X"A6",X"C8",X"5F",X"ED",X"C8",X"32",X"6F",X"C8",X"4A",X"A6",X"C8",X"53",X"26",
		X"08",X"EC",X"C8",X"34",X"E3",X"C8",X"30",X"20",X"20",X"EC",X"C8",X"34",X"2D",X"0C",X"27",X"1C",
		X"E3",X"C8",X"30",X"A1",X"C8",X"5E",X"22",X"0E",X"20",X"0F",X"E3",X"C8",X"30",X"A1",X"C8",X"5E",
		X"25",X"04",X"81",X"F0",X"25",X"03",X"A6",X"C8",X"5E",X"ED",X"C8",X"30",X"7E",X"1A",X"20",X"8E",
		X"1A",X"12",X"AF",X"C8",X"3E",X"96",X"39",X"27",X"09",X"A7",X"C8",X"44",X"CC",X"1A",X"27",X"7E",
		X"19",X"B4",X"A6",X"C8",X"58",X"27",X"0D",X"A6",X"C8",X"42",X"8E",X"1A",X"21",X"AE",X"86",X"AF",
		X"42",X"7E",X"19",X"E3",X"EC",X"C8",X"34",X"2D",X"2B",X"2E",X"07",X"63",X"C8",X"3A",X"2D",X"33",
		X"2A",X"0F",X"A6",X"C8",X"44",X"27",X"0A",X"6F",X"C8",X"44",X"86",X"04",X"A7",X"C8",X"45",X"20",
		X"36",X"A6",X"C8",X"45",X"8B",X"FE",X"2A",X"02",X"86",X"04",X"A7",X"C8",X"45",X"8E",X"1A",X"2D",
		X"EC",X"86",X"20",X"20",X"A6",X"C8",X"44",X"27",X"0A",X"6F",X"C8",X"44",X"86",X"04",X"A7",X"C8",
		X"45",X"20",X"14",X"A6",X"C8",X"45",X"8B",X"FE",X"2A",X"02",X"86",X"04",X"A7",X"C8",X"45",X"8E",
		X"1A",X"45",X"EC",X"86",X"ED",X"C8",X"40",X"A6",X"C8",X"32",X"81",X"A0",X"22",X"09",X"81",X"58",
		X"22",X"0A",X"CC",X"04",X"04",X"20",X"08",X"CC",X"00",X"00",X"20",X"03",X"CC",X"02",X"00",X"A7",
		X"C8",X"42",X"E7",X"C8",X"2A",X"8E",X"1A",X"5D",X"AE",X"86",X"AF",X"46",X"AE",X"C8",X"40",X"AE",
		X"86",X"AF",X"42",X"A6",X"46",X"44",X"40",X"AB",X"C8",X"30",X"A7",X"44",X"86",X"2A",X"E6",X"C8",
		X"31",X"2D",X"02",X"86",X"0A",X"A7",X"40",X"A6",X"47",X"44",X"40",X"AB",X"C8",X"32",X"A7",X"45",
		X"6C",X"4F",X"A6",X"C8",X"56",X"2A",X"19",X"AE",X"C8",X"54",X"A6",X"C8",X"42",X"A7",X"88",X"3B",
		X"20",X"0E",X"6A",X"C8",X"3B",X"2A",X"09",X"A6",X"C8",X"3C",X"A7",X"C8",X"3B",X"7E",X"14",X"8F",
		X"39",X"0C",X"A0",X"14",X"13",X"19",X"E5",X"07",X"FC",X"10",X"7B",X"17",X"15",X"1A",X"3F",X"1A",
		X"39",X"1A",X"33",X"09",X"25",X"11",X"61",X"17",X"C9",X"0A",X"4E",X"12",X"47",X"18",X"7D",X"0B",
		X"77",X"13",X"2D",X"19",X"31",X"1A",X"57",X"1A",X"51",X"1A",X"4B",X"04",X"81",X"0D",X"C9",X"14",
		X"F9",X"05",X"AA",X"0E",X"AF",X"15",X"AD",X"06",X"D3",X"0F",X"95",X"16",X"61",X"0B",X"1B",X"0A",
		X"17",X"09",X"14",X"16",X"A4",X"16",X"AE",X"16",X"B7",X"16",X"C0",X"16",X"C9",X"16",X"D2",X"16",
		X"DD",X"16",X"E8",X"16",X"F3",X"17",X"A3",X"17",X"A3",X"17",X"41",X"17",X"59",X"17",X"A7",X"17",
		X"A7",X"17",X"50",X"17",X"68",X"17",X"AB",X"18",X"3C",X"18",X"44",X"17",X"BB",X"17",X"CB",X"17",
		X"C3",X"18",X"2C",X"18",X"34",X"17",X"B3",X"17",X"D3",X"17",X"FC",X"18",X"04",X"18",X"78",X"18",
		X"8C",X"08",X"6C",X"5F",X"13",X"05",X"16",X"17",X"85",X"08",X"21",X"5E",X"A5",X"05",X"16",X"17",
		X"85",X"08",X"6B",X"5F",X"13",X"05",X"16",X"17",X"85",X"08",X"23",X"5E",X"A5",X"05",X"16",X"17",
		X"85",X"14",X"21",X"04",X"81",X"01",X"01",X"18",X"9E",X"10",X"00",X"41",X"8B",X"05",X"10",X"17",
		X"0F",X"10",X"00",X"41",X"DB",X"05",X"10",X"17",X"85",X"10",X"10",X"42",X"2B",X"07",X"19",X"17",
		X"19",X"10",X"10",X"42",X"DA",X"07",X"19",X"17",X"23",X"10",X"10",X"43",X"89",X"07",X"19",X"17",
		X"85",X"10",X"7D",X"44",X"38",X"07",X"19",X"17",X"2D",X"10",X"7D",X"44",X"E7",X"07",X"19",X"17",
		X"37",X"10",X"7D",X"45",X"96",X"07",X"19",X"17",X"85",X"10",X"31",X"00",X"2D",X"06",X"10",X"17",
		X"8F",X"10",X"32",X"00",X"8D",X"06",X"10",X"17",X"85",X"10",X"5C",X"00",X"2D",X"06",X"10",X"17",
		X"99",X"10",X"5B",X"00",X"8D",X"06",X"10",X"17",X"85",X"F0",X"00",X"F6",X"00",X"FA",X"00",X"FD",
		X"00",X"00",X"40",X"03",X"00",X"06",X"00",X"0A",X"00",X"10",X"00",X"00",X"00",X"F8",X"00",X"FB",
		X"00",X"FD",X"00",X"FE",X"80",X"00",X"40",X"01",X"80",X"03",X"00",X"05",X"00",X"08",X"00",X"00",
		X"00",X"39",X"86",X"01",X"A7",X"C8",X"1F",X"CC",X"1F",X"73",X"ED",X"C8",X"40",X"CC",X"00",X"00",
		X"A7",X"4E",X"A7",X"C8",X"1D",X"ED",X"C8",X"34",X"ED",X"C8",X"36",X"A7",X"C8",X"38",X"A7",X"C8",
		X"43",X"A7",X"C8",X"44",X"A7",X"C8",X"45",X"A7",X"C8",X"4A",X"A7",X"C8",X"4B",X"ED",X"C8",X"4C",
		X"A7",X"C8",X"4E",X"B6",X"A8",X"D9",X"A7",X"C8",X"3C",X"A7",X"C8",X"3B",X"8E",X"1B",X"AB",X"AF",
		X"C8",X"3E",X"8E",X"1B",X"98",X"AF",X"4A",X"39",X"A6",X"4E",X"27",X"04",X"BD",X"30",X"7C",X"39",
		X"A6",X"C8",X"4E",X"27",X"03",X"7E",X"1F",X"4C",X"6E",X"D8",X"3E",X"A6",X"C8",X"4B",X"27",X"03",
		X"7E",X"1F",X"1D",X"8E",X"1C",X"2A",X"AF",X"C8",X"3E",X"EC",X"C8",X"14",X"ED",X"C8",X"5E",X"E1",
		X"C8",X"32",X"25",X"1D",X"22",X"21",X"10",X"8E",X"00",X"00",X"A1",X"C8",X"30",X"26",X"1C",X"A6",
		X"C8",X"1D",X"26",X"53",X"86",X"FF",X"A7",X"C8",X"1D",X"BD",X"39",X"13",X"8E",X"00",X"00",X"20",
		X"3F",X"10",X"BE",X"A8",X"D7",X"20",X"04",X"10",X"BE",X"A8",X"D5",X"E6",X"C8",X"43",X"27",X"06",
		X"5A",X"E7",X"C8",X"43",X"20",X"10",X"9E",X"D5",X"8C",X"F4",X"00",X"23",X"12",X"0D",X"96",X"26",
		X"0E",X"C6",X"04",X"E7",X"C8",X"43",X"8E",X"00",X"00",X"10",X"8E",X"00",X"00",X"20",X"11",X"A1",
		X"C8",X"30",X"25",X"04",X"22",X"07",X"20",X"B7",X"BE",X"A8",X"D7",X"20",X"03",X"BE",X"A8",X"D5",
		X"10",X"AF",X"C8",X"36",X"AF",X"C8",X"34",X"7E",X"1F",X"1C",X"8E",X"1D",X"6F",X"AF",X"C8",X"3E",
		X"A6",X"C8",X"30",X"E6",X"C8",X"32",X"BD",X"67",X"5E",X"A7",X"C8",X"38",X"27",X"08",X"A7",X"C8",
		X"16",X"8E",X"1C",X"49",X"AF",X"4A",X"7E",X"1F",X"1C",X"A6",X"C8",X"16",X"8E",X"1F",X"B1",X"AE",
		X"86",X"A6",X"C8",X"30",X"E6",X"C8",X"32",X"6E",X"84",X"10",X"A3",X"C8",X"5E",X"27",X"08",X"20",
		X"23",X"10",X"A3",X"C8",X"5E",X"26",X"25",X"AE",X"C8",X"4C",X"27",X"0C",X"CC",X"00",X"00",X"A7",
		X"88",X"4B",X"A7",X"88",X"4E",X"ED",X"88",X"4C",X"BD",X"F9",X"16",X"39",X"C1",X"EC",X"25",X"5D",
		X"C6",X"EC",X"20",X"3F",X"C1",X"B1",X"22",X"55",X"C6",X"B1",X"20",X"27",X"C1",X"39",X"25",X"04",
		X"C6",X"39",X"20",X"2F",X"C1",X"37",X"22",X"45",X"C6",X"37",X"20",X"17",X"C1",X"38",X"22",X"3D",
		X"C6",X"38",X"20",X"0F",X"C1",X"97",X"22",X"35",X"C6",X"98",X"8E",X"00",X"00",X"AF",X"C8",X"34",
		X"BD",X"39",X"2F",X"E7",X"C8",X"32",X"EC",X"C8",X"36",X"2A",X"22",X"CC",X"00",X"00",X"ED",X"C8",
		X"36",X"20",X"1A",X"E7",X"C8",X"32",X"EC",X"C8",X"36",X"2F",X"12",X"20",X"EE",X"C1",X"68",X"25",
		X"0C",X"C6",X"68",X"20",X"EE",X"C1",X"48",X"25",X"04",X"C6",X"48",X"20",X"E6",X"CC",X"1B",X"98",
		X"ED",X"4A",X"39",X"A7",X"C8",X"30",X"EC",X"C8",X"34",X"2A",X"F2",X"CC",X"00",X"00",X"ED",X"C8",
		X"34",X"20",X"EA",X"A7",X"C8",X"30",X"EC",X"C8",X"34",X"2F",X"E2",X"20",X"EE",X"81",X"23",X"22",
		X"DC",X"86",X"23",X"20",X"DE",X"81",X"71",X"25",X"D4",X"86",X"71",X"20",X"E6",X"81",X"1E",X"22",
		X"CC",X"86",X"1E",X"20",X"CE",X"81",X"75",X"25",X"C4",X"86",X"75",X"20",X"D6",X"81",X"25",X"22",
		X"BC",X"86",X"25",X"8D",X"3C",X"20",X"BC",X"81",X"6E",X"25",X"B2",X"86",X"6E",X"8D",X"32",X"20",
		X"C2",X"81",X"27",X"22",X"A8",X"86",X"27",X"8D",X"28",X"20",X"A8",X"81",X"6C",X"25",X"9E",X"86",
		X"6C",X"8D",X"1E",X"20",X"AE",X"C6",X"10",X"E7",X"C8",X"14",X"E6",X"C8",X"32",X"E7",X"C8",X"15",
		X"86",X"01",X"20",X"8F",X"C6",X"80",X"E7",X"C8",X"14",X"E6",X"C8",X"32",X"E7",X"C8",X"15",X"20",
		X"92",X"D6",X"38",X"27",X"09",X"EC",X"C8",X"14",X"A7",X"C8",X"30",X"E7",X"C8",X"32",X"39",X"8E",
		X"1D",X"D4",X"AF",X"C8",X"3E",X"EC",X"C8",X"36",X"2D",X"23",X"26",X"17",X"EC",X"C8",X"34",X"26",
		X"2A",X"6C",X"C8",X"4A",X"A6",X"C8",X"4A",X"81",X"08",X"25",X"46",X"BD",X"39",X"2F",X"6F",X"C8",
		X"4A",X"20",X"3E",X"E3",X"C8",X"32",X"A1",X"C8",X"5F",X"22",X"0A",X"20",X"0B",X"E3",X"C8",X"32",
		X"A1",X"C8",X"5F",X"24",X"03",X"A6",X"C8",X"5F",X"ED",X"C8",X"32",X"6F",X"C8",X"4A",X"EC",X"C8",
		X"34",X"2D",X"0C",X"27",X"1C",X"E3",X"C8",X"30",X"A1",X"C8",X"5E",X"22",X"0E",X"20",X"0F",X"E3",
		X"C8",X"30",X"A1",X"C8",X"5E",X"25",X"04",X"81",X"F0",X"25",X"03",X"A6",X"C8",X"5E",X"ED",X"C8",
		X"30",X"7E",X"1F",X"1C",X"8E",X"1E",X"7C",X"AF",X"C8",X"3E",X"EC",X"C8",X"34",X"BD",X"1E",X"27",
		X"A6",X"C8",X"32",X"81",X"A0",X"22",X"08",X"81",X"58",X"22",X"07",X"86",X"04",X"20",X"05",X"4F",
		X"20",X"02",X"86",X"02",X"AE",X"C8",X"40",X"AE",X"86",X"AF",X"42",X"8E",X"1F",X"AD",X"AE",X"86",
		X"AF",X"46",X"8D",X"05",X"6C",X"4F",X"7E",X"1F",X"1C",X"A6",X"46",X"44",X"40",X"AB",X"C8",X"30",
		X"A7",X"44",X"86",X"2A",X"E6",X"C8",X"31",X"2D",X"02",X"86",X"0A",X"A7",X"40",X"A6",X"47",X"44",
		X"40",X"AB",X"C8",X"32",X"A7",X"45",X"39",X"2D",X"2F",X"2E",X"0B",X"86",X"FF",X"A7",X"C8",X"44",
		X"CC",X"1F",X"73",X"7E",X"1E",X"78",X"A6",X"C8",X"44",X"27",X"0A",X"6F",X"C8",X"44",X"86",X"02",
		X"A7",X"C8",X"45",X"20",X"0C",X"A6",X"C8",X"45",X"8B",X"FE",X"2A",X"02",X"86",X"06",X"A7",X"C8",
		X"45",X"8E",X"1F",X"79",X"EC",X"86",X"20",X"20",X"A6",X"C8",X"44",X"27",X"0A",X"6F",X"C8",X"44",
		X"86",X"02",X"A7",X"C8",X"45",X"20",X"0C",X"A6",X"C8",X"45",X"8B",X"FE",X"2A",X"02",X"86",X"06",
		X"A7",X"C8",X"45",X"8E",X"1F",X"93",X"EC",X"86",X"ED",X"C8",X"40",X"39",X"8E",X"1F",X"0E",X"AF",
		X"C8",X"3E",X"DC",X"D5",X"10",X"93",X"D9",X"25",X"21",X"AE",X"C8",X"4C",X"26",X"1C",X"BE",X"B0",
		X"09",X"27",X"09",X"8D",X"5D",X"27",X"15",X"AE",X"88",X"1A",X"26",X"F7",X"BE",X"B0",X"0D",X"27",
		X"09",X"8D",X"4F",X"27",X"07",X"AE",X"88",X"1A",X"26",X"F7",X"20",X"70",X"A6",X"0E",X"26",X"FA",
		X"A6",X"88",X"4E",X"27",X"19",X"96",X"D5",X"81",X"3C",X"22",X"EF",X"CC",X"00",X"00",X"A7",X"88",
		X"4E",X"10",X"AE",X"88",X"4C",X"ED",X"A8",X"4C",X"A7",X"A8",X"4B",X"A7",X"A8",X"4E",X"A6",X"C8",
		X"30",X"E6",X"C8",X"32",X"ED",X"88",X"14",X"AF",X"C8",X"4C",X"86",X"04",X"A7",X"C8",X"43",X"86",
		X"FF",X"A7",X"88",X"1E",X"6F",X"88",X"1D",X"A7",X"88",X"4B",X"EF",X"88",X"4C",X"6F",X"88",X"2B",
		X"20",X"B8",X"A6",X"88",X"30",X"A0",X"C8",X"30",X"2A",X"01",X"40",X"81",X"08",X"22",X"0E",X"A6",
		X"88",X"32",X"A0",X"C8",X"32",X"2A",X"01",X"40",X"81",X"10",X"22",X"01",X"4F",X"39",X"6A",X"C8",
		X"3B",X"2A",X"09",X"A6",X"C8",X"3C",X"A7",X"C8",X"3B",X"7E",X"1B",X"AB",X"39",X"8E",X"1F",X"0E",
		X"AF",X"C8",X"3E",X"8D",X"04",X"6C",X"4F",X"20",X"F3",X"96",X"D5",X"81",X"C0",X"25",X"04",X"96",
		X"D6",X"20",X"01",X"4F",X"BD",X"1E",X"27",X"AE",X"C8",X"4C",X"A6",X"88",X"42",X"AE",X"C8",X"40",
		X"AE",X"86",X"AF",X"42",X"8E",X"1F",X"AD",X"AE",X"86",X"AF",X"46",X"39",X"6F",X"C8",X"4E",X"AE",
		X"C8",X"4C",X"A6",X"88",X"30",X"E6",X"88",X"34",X"2B",X"04",X"9B",X"EF",X"20",X"02",X"9B",X"EE",
		X"A7",X"C8",X"30",X"E6",X"88",X"32",X"CB",X"05",X"E7",X"C8",X"32",X"8D",X"BC",X"BD",X"1E",X"09",
		X"6C",X"4F",X"39",X"25",X"0D",X"2A",X"9F",X"1C",X"13",X"1F",X"87",X"1F",X"8D",X"1F",X"87",X"1F",
		X"81",X"20",X"2D",X"2B",X"39",X"1C",X"7F",X"20",X"FD",X"2B",X"D3",X"1C",X"EB",X"21",X"CD",X"2C",
		X"6D",X"1D",X"57",X"1F",X"A1",X"1F",X"A7",X"1F",X"A1",X"1F",X"9B",X"22",X"9D",X"28",X"D1",X"1A",
		X"CF",X"23",X"6D",X"29",X"6B",X"1B",X"3B",X"24",X"3D",X"2A",X"05",X"1B",X"A7",X"08",X"1A",X"07",
		X"16",X"06",X"12",X"1C",X"8C",X"1C",X"94",X"1C",X"9C",X"1C",X"94",X"1C",X"8C",X"1C",X"84",X"1C",
		X"84",X"1C",X"9C",X"1C",X"9C",X"1C",X"59",X"1C",X"59",X"1D",X"1D",X"1D",X"27",X"1C",X"61",X"1C",
		X"61",X"1D",X"31",X"1D",X"3B",X"1C",X"7C",X"1D",X"0D",X"1D",X"15",X"1C",X"8C",X"1C",X"9C",X"1C",
		X"94",X"1C",X"FD",X"1D",X"05",X"1C",X"84",X"1C",X"A4",X"1C",X"CD",X"1C",X"D5",X"1D",X"45",X"1D",
		X"54",X"86",X"01",X"A7",X"C8",X"1F",X"CC",X"23",X"95",X"ED",X"C8",X"40",X"CC",X"00",X"00",X"A7",
		X"4E",X"A7",X"C8",X"1D",X"ED",X"C8",X"34",X"ED",X"C8",X"36",X"A7",X"C8",X"38",X"A7",X"C8",X"43",
		X"A7",X"C8",X"44",X"A7",X"C8",X"45",X"A7",X"C8",X"49",X"A7",X"C8",X"46",X"A7",X"C8",X"4A",X"B6",
		X"A8",X"D9",X"A7",X"C8",X"3C",X"A7",X"C8",X"3B",X"8E",X"20",X"37",X"AF",X"C8",X"3E",X"8E",X"20",
		X"34",X"AF",X"4A",X"39",X"6E",X"D8",X"3E",X"A6",X"4E",X"27",X"07",X"6F",X"C8",X"16",X"BD",X"30",
		X"7C",X"39",X"8E",X"20",X"BD",X"A6",X"C8",X"49",X"27",X"03",X"8E",X"23",X"11",X"AF",X"C8",X"3E",
		X"EC",X"C8",X"14",X"ED",X"C8",X"5E",X"E1",X"C8",X"32",X"25",X"1D",X"22",X"21",X"10",X"8E",X"00",
		X"00",X"A1",X"C8",X"30",X"26",X"1C",X"A6",X"C8",X"1D",X"26",X"4F",X"86",X"FF",X"A7",X"C8",X"1D",
		X"BD",X"39",X"13",X"8E",X"00",X"00",X"20",X"3B",X"10",X"BE",X"A8",X"D7",X"20",X"04",X"10",X"BE",
		X"A8",X"D5",X"E6",X"C8",X"43",X"27",X"06",X"5A",X"E7",X"C8",X"43",X"20",X"0C",X"9E",X"D5",X"8C",
		X"F0",X"00",X"23",X"0E",X"C6",X"04",X"E7",X"C8",X"43",X"8E",X"00",X"00",X"10",X"8E",X"00",X"00",
		X"20",X"11",X"A1",X"C8",X"30",X"25",X"04",X"22",X"07",X"20",X"BB",X"BE",X"A8",X"D7",X"20",X"03",
		X"BE",X"A8",X"D5",X"10",X"AF",X"C8",X"36",X"AF",X"C8",X"34",X"7E",X"23",X"10",X"8E",X"21",X"FD",
		X"AF",X"C8",X"3E",X"96",X"E3",X"81",X"11",X"27",X"08",X"96",X"39",X"26",X"0A",X"96",X"DB",X"26",
		X"06",X"96",X"D2",X"27",X"10",X"0F",X"D2",X"8E",X"70",X"A5",X"BD",X"6F",X"D3",X"86",X"FF",X"A7",
		X"C8",X"49",X"7E",X"23",X"10",X"A6",X"C8",X"30",X"E6",X"C8",X"32",X"BD",X"67",X"5E",X"A7",X"C8",
		X"38",X"27",X"08",X"A7",X"C8",X"16",X"8E",X"20",X"FE",X"AF",X"4A",X"7E",X"23",X"10",X"A6",X"C8",
		X"16",X"8E",X"23",X"F7",X"AE",X"86",X"A6",X"C8",X"30",X"E6",X"C8",X"32",X"6E",X"84",X"10",X"A3",
		X"C8",X"5E",X"27",X"08",X"20",X"12",X"10",X"A3",X"C8",X"5E",X"26",X"14",X"BD",X"F9",X"16",X"39",
		X"C1",X"EC",X"25",X"5D",X"C6",X"EC",X"20",X"3F",X"C1",X"B1",X"22",X"55",X"C6",X"B1",X"20",X"27",
		X"C1",X"39",X"25",X"04",X"C6",X"39",X"20",X"2F",X"C1",X"37",X"22",X"45",X"C6",X"37",X"20",X"17",
		X"C1",X"38",X"22",X"3D",X"C6",X"38",X"20",X"0F",X"C1",X"97",X"22",X"35",X"C6",X"98",X"8E",X"00",
		X"00",X"AF",X"C8",X"34",X"BD",X"39",X"2F",X"E7",X"C8",X"32",X"EC",X"C8",X"36",X"2A",X"22",X"CC",
		X"00",X"00",X"ED",X"C8",X"36",X"20",X"1A",X"E7",X"C8",X"32",X"EC",X"C8",X"36",X"2F",X"12",X"20",
		X"EE",X"C1",X"68",X"25",X"0C",X"C6",X"68",X"20",X"EE",X"C1",X"48",X"25",X"04",X"C6",X"48",X"20",
		X"E6",X"CC",X"20",X"34",X"ED",X"4A",X"39",X"A7",X"C8",X"30",X"EC",X"C8",X"34",X"2A",X"F2",X"CC",
		X"00",X"00",X"ED",X"C8",X"34",X"20",X"EA",X"A7",X"C8",X"30",X"EC",X"C8",X"34",X"2F",X"E2",X"20",
		X"EE",X"81",X"23",X"22",X"DC",X"86",X"23",X"20",X"DE",X"81",X"6F",X"25",X"D4",X"86",X"6F",X"20",
		X"E6",X"81",X"1E",X"22",X"CC",X"86",X"1E",X"20",X"CE",X"81",X"75",X"25",X"C4",X"86",X"75",X"20",
		X"D6",X"81",X"25",X"22",X"BC",X"86",X"25",X"20",X"BE",X"81",X"6E",X"25",X"B4",X"86",X"6E",X"20",
		X"C6",X"81",X"27",X"22",X"AC",X"86",X"27",X"20",X"AE",X"81",X"6C",X"25",X"A4",X"86",X"6C",X"20",
		X"B6",X"C6",X"10",X"E7",X"C8",X"14",X"E6",X"C8",X"32",X"E7",X"C8",X"15",X"86",X"01",X"20",X"97",
		X"C6",X"80",X"E7",X"C8",X"14",X"E6",X"C8",X"32",X"E7",X"C8",X"15",X"20",X"9A",X"8E",X"22",X"5F",
		X"AF",X"C8",X"3E",X"EC",X"C8",X"36",X"2D",X"20",X"26",X"14",X"EC",X"C8",X"34",X"26",X"27",X"6C",
		X"C8",X"4A",X"A6",X"C8",X"4A",X"81",X"08",X"25",X"43",X"BD",X"39",X"2F",X"20",X"3E",X"E3",X"C8",
		X"32",X"A1",X"C8",X"5F",X"22",X"0A",X"20",X"0B",X"E3",X"C8",X"32",X"A1",X"C8",X"5F",X"24",X"03",
		X"A6",X"C8",X"5F",X"ED",X"C8",X"32",X"6F",X"C8",X"4A",X"EC",X"C8",X"34",X"2D",X"0C",X"27",X"1C",
		X"E3",X"C8",X"30",X"A1",X"C8",X"5E",X"22",X"0E",X"20",X"0F",X"E3",X"C8",X"30",X"A1",X"C8",X"5E",
		X"25",X"04",X"81",X"F0",X"25",X"03",X"A6",X"C8",X"5E",X"ED",X"C8",X"30",X"7E",X"23",X"10",X"8E",
		X"23",X"02",X"AF",X"C8",X"3E",X"EC",X"C8",X"34",X"2D",X"2F",X"2E",X"0B",X"86",X"FF",X"A7",X"C8",
		X"44",X"CC",X"23",X"95",X"7E",X"22",X"B9",X"A6",X"C8",X"44",X"27",X"0A",X"6F",X"C8",X"44",X"86",
		X"02",X"A7",X"C8",X"45",X"20",X"0C",X"A6",X"C8",X"45",X"8B",X"FE",X"2A",X"02",X"86",X"06",X"A7",
		X"C8",X"45",X"8E",X"23",X"9B",X"EC",X"86",X"20",X"20",X"A6",X"C8",X"44",X"27",X"0A",X"6F",X"C8",
		X"44",X"86",X"02",X"A7",X"C8",X"45",X"20",X"0C",X"A6",X"C8",X"45",X"8B",X"FE",X"2A",X"02",X"86",
		X"06",X"A7",X"C8",X"45",X"8E",X"23",X"B5",X"EC",X"86",X"ED",X"C8",X"40",X"8D",X"2F",X"AE",X"C8",
		X"40",X"AE",X"86",X"AF",X"42",X"8E",X"23",X"CF",X"AE",X"86",X"AF",X"46",X"A6",X"46",X"44",X"40",
		X"AB",X"C8",X"30",X"A7",X"44",X"86",X"2A",X"E6",X"C8",X"31",X"2D",X"02",X"86",X"0A",X"A7",X"40",
		X"A6",X"47",X"44",X"40",X"AB",X"C8",X"32",X"A7",X"45",X"6C",X"4F",X"20",X"23",X"A6",X"C8",X"32",
		X"81",X"A0",X"22",X"08",X"81",X"58",X"22",X"07",X"86",X"04",X"20",X"05",X"4F",X"20",X"02",X"86",
		X"02",X"39",X"6A",X"C8",X"3B",X"2A",X"09",X"A6",X"C8",X"3C",X"A7",X"C8",X"3B",X"7E",X"20",X"37",
		X"39",X"8E",X"23",X"02",X"AF",X"C8",X"3E",X"8E",X"23",X"23",X"A6",X"C8",X"46",X"48",X"AD",X"96",
		X"7E",X"23",X"10",X"23",X"31",X"23",X"38",X"23",X"3D",X"23",X"46",X"23",X"4F",X"23",X"58",X"23",
		X"94",X"86",X"00",X"A7",X"C8",X"3C",X"20",X"59",X"8E",X"23",X"95",X"20",X"4B",X"8E",X"23",X"D5",
		X"10",X"8E",X"23",X"E7",X"20",X"37",X"8E",X"23",X"DB",X"10",X"8E",X"23",X"ED",X"20",X"2E",X"8E",
		X"23",X"E1",X"10",X"8E",X"23",X"F3",X"20",X"25",X"86",X"FF",X"A7",X"C8",X"16",X"BD",X"30",X"7C",
		X"10",X"8E",X"49",X"80",X"A6",X"C8",X"30",X"E6",X"C8",X"32",X"1F",X"01",X"4F",X"C6",X"04",X"34",
		X"40",X"BD",X"63",X"61",X"86",X"FF",X"A7",X"C8",X"1E",X"35",X"40",X"20",X"14",X"BD",X"22",X"ED",
		X"10",X"AE",X"A6",X"10",X"AF",X"46",X"20",X"03",X"BD",X"22",X"ED",X"AE",X"86",X"AF",X"42",X"6C",
		X"4F",X"6C",X"C8",X"46",X"39",X"25",X"0D",X"2A",X"9F",X"1C",X"13",X"23",X"A9",X"23",X"AF",X"23",
		X"A9",X"23",X"A3",X"20",X"2D",X"2B",X"39",X"1C",X"7F",X"20",X"FD",X"2B",X"D3",X"1C",X"EB",X"21",
		X"CD",X"2C",X"6D",X"1D",X"57",X"23",X"C3",X"23",X"C9",X"23",X"C3",X"23",X"BD",X"22",X"9D",X"28",
		X"D1",X"1A",X"CF",X"23",X"6D",X"29",X"6B",X"1B",X"3B",X"24",X"3D",X"2A",X"05",X"1B",X"A7",X"08",
		X"1A",X"07",X"16",X"06",X"12",X"25",X"DD",X"2D",X"07",X"1D",X"C3",X"26",X"D9",X"2D",X"E8",X"1E",
		X"63",X"27",X"D5",X"2E",X"C9",X"1F",X"03",X"09",X"1C",X"09",X"19",X"08",X"14",X"09",X"1C",X"09",
		X"19",X"08",X"14",X"09",X"1C",X"09",X"19",X"08",X"14",X"21",X"30",X"21",X"38",X"21",X"40",X"21",
		X"38",X"21",X"30",X"21",X"28",X"21",X"28",X"21",X"40",X"21",X"40",X"21",X"0E",X"21",X"0E",X"21",
		X"C1",X"21",X"C9",X"21",X"16",X"21",X"16",X"21",X"D1",X"21",X"D9",X"21",X"20",X"21",X"B1",X"21",
		X"B9",X"21",X"30",X"21",X"40",X"21",X"38",X"21",X"A1",X"21",X"A9",X"21",X"28",X"21",X"48",X"21",
		X"71",X"21",X"79",X"21",X"E1",X"21",X"F0",X"8E",X"26",X"D7",X"86",X"05",X"8D",X"51",X"CC",X"00",
		X"00",X"ED",X"C8",X"4D",X"39",X"8E",X"26",X"C0",X"86",X"01",X"8D",X"43",X"CC",X"20",X"0B",X"8E",
		X"72",X"5E",X"8D",X"11",X"39",X"8E",X"26",X"EE",X"86",X"01",X"8D",X"33",X"CC",X"23",X"0E",X"8E",
		X"6E",X"5A",X"8D",X"01",X"39",X"ED",X"C8",X"3D",X"AF",X"C8",X"3F",X"30",X"C4",X"34",X"40",X"BD",
		X"F8",X"B5",X"86",X"24",X"A7",X"4C",X"CC",X"12",X"00",X"ED",X"40",X"A6",X"05",X"4C",X"A7",X"45",
		X"CC",X"01",X"01",X"ED",X"46",X"EF",X"88",X"4D",X"CC",X"24",X"64",X"ED",X"4A",X"35",X"C0",X"A7",
		X"C8",X"1F",X"A6",X"00",X"5F",X"ED",X"40",X"E7",X"C8",X"4C",X"EC",X"03",X"ED",X"C8",X"3B",X"54",
		X"44",X"ED",X"C8",X"36",X"EC",X"01",X"ED",X"4A",X"ED",X"C8",X"41",X"EC",X"05",X"ED",X"C8",X"39",
		X"E6",X"C8",X"14",X"CB",X"20",X"E7",X"C8",X"38",X"E6",X"C8",X"30",X"CB",X"20",X"E1",X"C8",X"38",
		X"25",X"02",X"30",X"08",X"EC",X"07",X"ED",X"C8",X"34",X"EC",X"09",X"ED",X"C8",X"46",X"EC",X"0B",
		X"ED",X"C8",X"48",X"EC",X"0D",X"ED",X"C8",X"4A",X"6F",X"C8",X"43",X"A6",X"C8",X"32",X"A0",X"C8",
		X"37",X"A7",X"45",X"39",X"BD",X"26",X"98",X"BD",X"26",X"62",X"10",X"26",X"00",X"A8",X"BD",X"25",
		X"75",X"26",X"01",X"39",X"8E",X"70",X"C5",X"BD",X"6F",X"D3",X"8E",X"25",X"00",X"AF",X"4A",X"39",
		X"A6",X"C8",X"1D",X"27",X"09",X"BD",X"26",X"98",X"EC",X"C8",X"44",X"ED",X"42",X"39",X"AE",X"C8",
		X"41",X"AF",X"4A",X"8E",X"70",X"BD",X"BD",X"6F",X"D3",X"39",X"BD",X"26",X"98",X"BD",X"26",X"62",
		X"27",X"1B",X"7E",X"25",X"96",X"BD",X"26",X"98",X"BD",X"26",X"62",X"27",X"10",X"A6",X"C8",X"30",
		X"A0",X"C8",X"36",X"A7",X"44",X"EC",X"C8",X"3B",X"ED",X"46",X"7E",X"25",X"E4",X"BD",X"25",X"75",
		X"26",X"01",X"39",X"8E",X"70",X"C5",X"BD",X"6F",X"D3",X"8E",X"27",X"16",X"AF",X"C8",X"39",X"8E",
		X"25",X"55",X"AF",X"4A",X"39",X"A6",X"C8",X"1D",X"27",X"09",X"BD",X"26",X"98",X"EC",X"C8",X"44",
		X"ED",X"42",X"39",X"8E",X"27",X"0F",X"AF",X"C8",X"39",X"AE",X"C8",X"41",X"AF",X"4A",X"8E",X"70",
		X"BD",X"BD",X"6F",X"D3",X"39",X"86",X"FF",X"A7",X"C8",X"1D",X"EC",X"C8",X"14",X"81",X"AD",X"25",
		X"14",X"81",X"F2",X"22",X"10",X"AD",X"D8",X"22",X"34",X"40",X"EE",X"C8",X"4D",X"27",X"03",X"BD",
		X"F9",X"4B",X"35",X"40",X"4F",X"39",X"EC",X"C8",X"30",X"A0",X"C8",X"36",X"A7",X"44",X"0D",X"E4",
		X"26",X"35",X"81",X"40",X"22",X"1B",X"A1",X"C8",X"3D",X"24",X"2C",X"A1",X"C8",X"3E",X"23",X"20",
		X"E6",X"C8",X"3E",X"AE",X"C8",X"4D",X"E7",X"04",X"EC",X"C8",X"3B",X"ED",X"06",X"ED",X"46",X"20",
		X"23",X"A1",X"C8",X"40",X"23",X"11",X"A1",X"C8",X"3F",X"22",X"05",X"E6",X"C8",X"3F",X"20",X"E3",
		X"CC",X"01",X"01",X"ED",X"46",X"20",X"05",X"EC",X"C8",X"3B",X"ED",X"46",X"AE",X"C8",X"4D",X"CC",
		X"01",X"01",X"ED",X"06",X"EC",X"C8",X"44",X"ED",X"42",X"A6",X"40",X"84",X"DF",X"6D",X"C8",X"31",
		X"2A",X"02",X"8A",X"20",X"A7",X"40",X"6C",X"4F",X"39",X"34",X"42",X"8D",X"26",X"27",X"07",X"8D",
		X"12",X"86",X"FF",X"A7",X"C8",X"4C",X"35",X"C2",X"EC",X"C8",X"34",X"58",X"49",X"ED",X"C8",X"34",
		X"8D",X"01",X"39",X"86",X"AD",X"6D",X"C8",X"34",X"2A",X"02",X"86",X"F2",X"A7",X"C8",X"14",X"6F",
		X"C8",X"1D",X"39",X"FE",X"B0",X"35",X"26",X"03",X"FE",X"B0",X"39",X"39",X"34",X"40",X"8D",X"F3",
		X"27",X"1B",X"CC",X"27",X"20",X"ED",X"C8",X"39",X"A6",X"C8",X"3B",X"E6",X"C8",X"34",X"2A",X"01",
		X"40",X"AB",X"C8",X"30",X"A7",X"C8",X"14",X"E6",X"C8",X"15",X"6F",X"C8",X"1D",X"35",X"C0",X"34",
		X"40",X"8D",X"D0",X"27",X"0B",X"A6",X"C8",X"34",X"97",X"98",X"A6",X"C8",X"30",X"E6",X"C8",X"32",
		X"35",X"C0",X"96",X"39",X"A4",X"C8",X"4C",X"26",X"12",X"EC",X"C8",X"34",X"2B",X"07",X"8D",X"0C",
		X"25",X"09",X"8D",X"1A",X"39",X"8D",X"05",X"22",X"02",X"8D",X"13",X"39",X"E3",X"C8",X"30",X"ED",
		X"C8",X"30",X"8B",X"1E",X"E6",X"C8",X"14",X"CB",X"1E",X"34",X"04",X"A1",X"E0",X"39",X"A6",X"C8",
		X"14",X"A7",X"C8",X"30",X"6F",X"C8",X"31",X"39",X"6A",X"C8",X"43",X"2E",X"22",X"AE",X"C8",X"39",
		X"EC",X"81",X"26",X"04",X"AE",X"84",X"EC",X"81",X"A7",X"C8",X"43",X"EB",X"C8",X"32",X"E0",X"C8",
		X"37",X"E7",X"45",X"E6",X"80",X"AF",X"C8",X"39",X"AE",X"C5",X"AF",X"C8",X"44",X"6C",X"4F",X"39",
		X"0A",X"25",X"1A",X"15",X"14",X"27",X"0F",X"01",X"00",X"5B",X"5D",X"5D",X"01",X"00",X"00",X"FF",
		X"00",X"58",X"15",X"59",X"B9",X"00",X"00",X"0A",X"25",X"25",X"18",X"17",X"27",X"0F",X"00",X"C0",
		X"0B",X"41",X"0D",X"69",X"00",X"00",X"FF",X"40",X"0F",X"91",X"11",X"B9",X"00",X"00",X"0A",X"24",
		X"E4",X"15",X"12",X"27",X"05",X"01",X"00",X"36",X"3A",X"37",X"B4",X"00",X"00",X"FF",X"00",X"33",
		X"46",X"34",X"C0",X"00",X"00",X"04",X"00",X"46",X"04",X"00",X"48",X"00",X"00",X"27",X"05",X"06",
		X"00",X"48",X"00",X"00",X"27",X"0F",X"05",X"00",X"46",X"05",X"00",X"48",X"00",X"00",X"27",X"16",
		X"02",X"00",X"46",X"00",X"00",X"27",X"20",X"34",X"66",X"BD",X"F3",X"66",X"27",X"05",X"8E",X"CD",
		X"00",X"20",X"03",X"8E",X"CC",X"00",X"34",X"10",X"10",X"8E",X"CD",X"FF",X"C6",X"05",X"BD",X"7F",
		X"26",X"AE",X"E4",X"A6",X"80",X"84",X"0F",X"81",X"05",X"26",X"20",X"8C",X"CE",X"00",X"25",X"F3",
		X"AE",X"E4",X"C6",X"0A",X"BD",X"7F",X"26",X"AE",X"E1",X"A6",X"80",X"84",X"0F",X"81",X"0A",X"26",
		X"0A",X"8C",X"CE",X"00",X"25",X"F3",X"8E",X"00",X"00",X"20",X"02",X"30",X"1F",X"35",X"E6",X"34",
		X"76",X"DE",X"AC",X"27",X"07",X"AD",X"D8",X"02",X"EE",X"44",X"26",X"F9",X"35",X"F6",X"DE",X"AC",
		X"27",X"06",X"6C",X"4F",X"EE",X"44",X"26",X"FA",X"BD",X"E5",X"1F",X"DC",X"AC",X"26",X"F9",X"39",
		X"DE",X"AC",X"27",X"06",X"8D",X"3A",X"EE",X"44",X"26",X"FA",X"39",X"34",X"31",X"1A",X"50",X"34",
		X"10",X"BE",X"AD",X"85",X"EE",X"81",X"26",X"07",X"35",X"10",X"35",X"31",X"86",X"FF",X"39",X"BF",
		X"AD",X"85",X"35",X"10",X"AF",X"42",X"10",X"AF",X"4A",X"6F",X"4E",X"6F",X"4F",X"CC",X"00",X"00",
		X"ED",X"46",X"9E",X"AC",X"DF",X"AC",X"AF",X"44",X"27",X"02",X"EF",X"06",X"35",X"31",X"4F",X"39",
		X"34",X"01",X"1A",X"50",X"BE",X"AD",X"85",X"EF",X"83",X"BF",X"AD",X"85",X"AE",X"46",X"26",X"0C",
		X"10",X"AE",X"44",X"10",X"9F",X"AC",X"27",X"02",X"AF",X"26",X"35",X"81",X"10",X"AE",X"44",X"10",
		X"AF",X"04",X"27",X"02",X"AF",X"26",X"35",X"81",X"34",X"57",X"1A",X"50",X"CE",X"AD",X"87",X"EF",
		X"5E",X"8E",X"AA",X"65",X"86",X"32",X"AF",X"C1",X"30",X"88",X"10",X"4A",X"26",X"F8",X"CC",X"00",
		X"00",X"ED",X"C4",X"DD",X"AC",X"35",X"D7",X"6F",X"4D",X"20",X"02",X"8D",X"0B",X"86",X"02",X"A7",
		X"C8",X"1E",X"CC",X"28",X"32",X"ED",X"4A",X"39",X"BD",X"3E",X"78",X"96",X"D5",X"84",X"1F",X"A7",
		X"4D",X"39",X"6A",X"4D",X"2E",X"11",X"6C",X"45",X"6A",X"47",X"26",X"04",X"AD",X"D8",X"22",X"39",
		X"A6",X"C8",X"1E",X"A7",X"4D",X"6C",X"4F",X"39",X"8D",X"DE",X"86",X"02",X"A7",X"C8",X"1E",X"A6",
		X"47",X"A7",X"C8",X"1D",X"6F",X"47",X"AB",X"45",X"A7",X"45",X"EC",X"4A",X"ED",X"C8",X"28",X"CC",
		X"28",X"65",X"ED",X"4A",X"39",X"6A",X"4D",X"2E",X"18",X"6A",X"45",X"6C",X"47",X"6A",X"C8",X"1D",
		X"26",X"08",X"AE",X"C8",X"28",X"AF",X"4A",X"6C",X"4F",X"39",X"A6",X"C8",X"1E",X"A7",X"4D",X"6C",
		X"4F",X"39",X"86",X"FF",X"A7",X"C8",X"46",X"CC",X"28",X"95",X"ED",X"C8",X"47",X"A6",X"40",X"8A",
		X"18",X"A7",X"40",X"20",X"18",X"6A",X"C8",X"45",X"2E",X"31",X"AE",X"C8",X"43",X"EC",X"81",X"26",
		X"22",X"6A",X"C8",X"40",X"27",X"07",X"AE",X"C8",X"41",X"EC",X"81",X"20",X"16",X"A6",X"80",X"26",
		X"0A",X"6F",X"C8",X"46",X"8E",X"28",X"CB",X"AF",X"C8",X"47",X"39",X"A7",X"C8",X"40",X"AF",X"C8",
		X"41",X"EC",X"81",X"E7",X"41",X"A7",X"C8",X"45",X"AF",X"C8",X"43",X"39",X"86",X"FF",X"A7",X"C8",
		X"56",X"CC",X"28",X"DE",X"ED",X"C8",X"57",X"EC",X"44",X"ED",X"C8",X"59",X"20",X"18",X"6A",X"C8",
		X"55",X"2E",X"3A",X"AE",X"C8",X"53",X"A6",X"80",X"26",X"22",X"6A",X"C8",X"50",X"27",X"07",X"AE",
		X"C8",X"51",X"A6",X"80",X"20",X"16",X"A6",X"80",X"26",X"0A",X"6F",X"C8",X"56",X"8E",X"29",X"1D",
		X"AF",X"C8",X"57",X"39",X"A7",X"C8",X"50",X"AF",X"C8",X"51",X"A6",X"80",X"A7",X"C8",X"55",X"EC",
		X"C8",X"59",X"AB",X"80",X"E0",X"80",X"ED",X"44",X"AF",X"C8",X"53",X"6C",X"4F",X"39",X"86",X"FF",
		X"97",X"F4",X"97",X"96",X"BD",X"2A",X"8A",X"BD",X"2A",X"AD",X"86",X"04",X"B7",X"BB",X"B7",X"B7",
		X"A8",X"F2",X"B7",X"AF",X"7E",X"B7",X"A8",X"F8",X"7F",X"A8",X"D9",X"BD",X"E5",X"1F",X"8E",X"2A",
		X"D6",X"BD",X"F5",X"CC",X"CC",X"00",X"3C",X"BD",X"2A",X"86",X"8E",X"2B",X"21",X"BD",X"F5",X"CC",
		X"86",X"3C",X"CE",X"2B",X"73",X"BD",X"2A",X"6B",X"BD",X"29",X"E3",X"BD",X"2A",X"8A",X"BD",X"2A",
		X"03",X"8E",X"2B",X"40",X"BD",X"F5",X"CC",X"CC",X"3E",X"06",X"BD",X"2A",X"59",X"86",X"FF",X"97",
		X"39",X"BD",X"29",X"E3",X"BD",X"2A",X"03",X"BD",X"2A",X"8A",X"86",X"14",X"CE",X"2B",X"97",X"BD",
		X"2A",X"7D",X"CE",X"2B",X"9D",X"BD",X"2A",X"75",X"CE",X"2B",X"A3",X"BD",X"2A",X"7D",X"CE",X"2B",
		X"A9",X"BD",X"2A",X"75",X"CE",X"2B",X"AF",X"BD",X"2A",X"7D",X"CE",X"2B",X"B5",X"BD",X"2A",X"7D",
		X"86",X"1E",X"BD",X"2A",X"A6",X"86",X"FF",X"97",X"39",X"97",X"E4",X"BD",X"00",X"B5",X"BD",X"29",
		X"E3",X"0F",X"39",X"CC",X"2D",X"08",X"BD",X"2A",X"59",X"BD",X"29",X"E3",X"BD",X"2A",X"03",X"CC",
		X"3E",X"04",X"BD",X"2A",X"59",X"86",X"FF",X"97",X"39",X"BD",X"29",X"E3",X"BD",X"2A",X"03",X"8E",
		X"2B",X"5E",X"BD",X"F5",X"CC",X"CC",X"00",X"B4",X"BD",X"2A",X"86",X"BD",X"00",X"B5",X"0F",X"E4",
		X"0F",X"F4",X"39",X"8D",X"19",X"C6",X"0C",X"34",X"04",X"8E",X"70",X"85",X"BD",X"6F",X"D3",X"96",
		X"D5",X"84",X"0F",X"8B",X"07",X"BD",X"2A",X"A6",X"6A",X"E4",X"26",X"ED",X"35",X"84",X"C6",X"FF",
		X"D7",X"9A",X"39",X"BD",X"00",X"B5",X"0F",X"39",X"BE",X"B0",X"09",X"27",X"02",X"8D",X"3B",X"BE",
		X"B0",X"0D",X"27",X"02",X"8D",X"34",X"BE",X"B0",X"11",X"27",X"02",X"8D",X"2D",X"BE",X"B0",X"15",
		X"27",X"02",X"8D",X"26",X"BE",X"B0",X"1D",X"27",X"02",X"8D",X"1F",X"BE",X"B0",X"19",X"27",X"02",
		X"8D",X"18",X"BD",X"E5",X"1F",X"F6",X"B0",X"08",X"FB",X"B0",X"0C",X"FB",X"B0",X"10",X"FB",X"B0",
		X"14",X"FB",X"B0",X"18",X"FB",X"B0",X"1C",X"26",X"E9",X"39",X"FC",X"51",X"29",X"ED",X"88",X"14",
		X"6F",X"88",X"1D",X"AE",X"88",X"1A",X"26",X"F2",X"39",X"CE",X"AE",X"6E",X"E7",X"41",X"E7",X"47",
		X"E7",X"4D",X"E7",X"C8",X"13",X"E7",X"C8",X"19",X"E7",X"C8",X"1F",X"C6",X"06",X"8D",X"06",X"33",
		X"46",X"5A",X"26",X"F9",X"39",X"34",X"02",X"8D",X"04",X"8D",X"2B",X"35",X"82",X"34",X"46",X"37",
		X"36",X"BD",X"63",X"61",X"35",X"C6",X"8D",X"0C",X"8D",X"13",X"BD",X"E5",X"1F",X"8E",X"2B",X"6D",
		X"BD",X"F4",X"87",X"39",X"BD",X"E5",X"1F",X"7D",X"BC",X"2D",X"2A",X"F8",X"39",X"BD",X"E5",X"1F",
		X"83",X"00",X"01",X"26",X"F8",X"39",X"BD",X"E5",X"1F",X"4A",X"26",X"FA",X"39",X"CE",X"2B",X"73",
		X"10",X"8E",X"AE",X"6E",X"8E",X"00",X"24",X"BD",X"7F",X"33",X"CC",X"21",X"31",X"B7",X"AE",X"72",
		X"F7",X"AE",X"78",X"CC",X"41",X"51",X"B7",X"AE",X"7E",X"F7",X"AE",X"84",X"CC",X"61",X"71",X"B7",
		X"AE",X"8A",X"F7",X"AE",X"90",X"39",X"2A",X"DC",X"00",X"55",X"6C",X"44",X"54",X"68",X"65",X"20",
		X"54",X"75",X"72",X"6B",X"65",X"79",X"20",X"53",X"68",X"6F",X"6F",X"74",X"5C",X"63",X"68",X"61",
		X"72",X"61",X"63",X"74",X"65",X"72",X"73",X"20",X"77",X"6F",X"75",X"6C",X"64",X"20",X"6E",X"6F",
		X"77",X"5C",X"6C",X"69",X"6B",X"65",X"20",X"74",X"6F",X"20",X"74",X"68",X"61",X"6E",X"6B",X"20",
		X"79",X"6F",X"75",X"20",X"66",X"6F",X"72",X"5C",X"70",X"6C",X"61",X"79",X"69",X"6E",X"67",X"2E",
		X"FF",X"2B",X"27",X"00",X"4C",X"6C",X"44",X"54",X"68",X"65",X"20",X"67",X"6F",X"6F",X"64",X"20",
		X"67",X"75",X"79",X"73",X"20",X"74",X"68",X"61",X"6E",X"6B",X"20",X"79",X"6F",X"75",X"2E",X"FF",
		X"2B",X"46",X"00",X"4F",X"6C",X"44",X"54",X"68",X"65",X"20",X"62",X"61",X"64",X"20",X"67",X"75",
		X"79",X"73",X"20",X"74",X"68",X"61",X"6E",X"6B",X"20",X"79",X"6F",X"75",X"2E",X"FF",X"2B",X"64",
		X"00",X"7C",X"6C",X"44",X"54",X"48",X"45",X"20",X"45",X"4E",X"44",X"3F",X"FF",X"00",X"00",X"4D",
		X"60",X"4D",X"60",X"00",X"0A",X"8F",X"CC",X"2B",X"B8",X"00",X"0A",X"8F",X"CC",X"37",X"B8",X"00",
		X"0E",X"8F",X"CC",X"43",X"B8",X"00",X"0E",X"8F",X"CC",X"4F",X"B8",X"00",X"0C",X"8F",X"CC",X"5B",
		X"B8",X"00",X"0C",X"8F",X"CC",X"67",X"B8",X"00",X"02",X"40",X"00",X"47",X"0A",X"00",X"02",X"50",
		X"00",X"4B",X"0A",X"00",X"02",X"30",X"00",X"43",X"0A",X"00",X"02",X"60",X"00",X"4F",X"0A",X"00",
		X"02",X"20",X"00",X"3F",X"0A",X"00",X"02",X"70",X"00",X"53",X"0A",X"86",X"01",X"A7",X"C8",X"1F",
		X"BD",X"63",X"23",X"AF",X"C8",X"54",X"CC",X"2F",X"70",X"ED",X"C8",X"40",X"CC",X"00",X"00",X"A7",
		X"4E",X"ED",X"C8",X"47",X"A7",X"C8",X"1D",X"ED",X"C8",X"34",X"ED",X"C8",X"36",X"A7",X"C8",X"38",
		X"A7",X"C8",X"42",X"A7",X"C8",X"44",X"A7",X"C8",X"45",X"A7",X"C8",X"4A",X"A7",X"C8",X"46",X"ED",
		X"C8",X"4E",X"86",X"07",X"A7",X"C8",X"4D",X"B6",X"A8",X"F8",X"A7",X"C8",X"3C",X"A7",X"C8",X"3B",
		X"8E",X"2C",X"0F",X"AF",X"C8",X"3E",X"8E",X"2C",X"0C",X"AF",X"4A",X"39",X"6E",X"D8",X"3E",X"A6",
		X"4E",X"27",X"0C",X"AE",X"C8",X"4E",X"27",X"03",X"6A",X"88",X"4F",X"BD",X"30",X"7C",X"39",X"8E",
		X"2C",X"E7",X"AF",X"C8",X"3E",X"AE",X"C8",X"4E",X"27",X"2D",X"A6",X"0C",X"81",X"20",X"27",X"0C",
		X"A6",X"0E",X"27",X"08",X"CC",X"00",X"00",X"ED",X"C8",X"4E",X"20",X"28",X"96",X"D5",X"C6",X"08",
		X"3D",X"D6",X"D6",X"2B",X"01",X"40",X"AB",X"88",X"30",X"D6",X"D6",X"C4",X"01",X"EB",X"88",X"32",
		X"CB",X"03",X"ED",X"C8",X"14",X"20",X"10",X"6A",X"C8",X"4D",X"26",X"08",X"86",X"07",X"A7",X"C8",
		X"4D",X"BD",X"2C",X"AD",X"EC",X"C8",X"14",X"ED",X"C8",X"5E",X"A1",X"C8",X"30",X"25",X"19",X"22",
		X"1C",X"8E",X"00",X"00",X"E1",X"C8",X"32",X"26",X"17",X"A6",X"C8",X"1D",X"26",X"2C",X"86",X"FF",
		X"A7",X"C8",X"1D",X"BD",X"39",X"13",X"20",X"0F",X"BE",X"A8",X"F6",X"20",X"03",X"BE",X"A8",X"F4",
		X"E1",X"C8",X"32",X"25",X"07",X"22",X"0A",X"CC",X"00",X"00",X"20",X"08",X"FC",X"A8",X"F6",X"20",
		X"03",X"FC",X"A8",X"F4",X"ED",X"C8",X"36",X"AF",X"C8",X"34",X"7E",X"2F",X"69",X"BE",X"B0",X"0D",
		X"27",X"0C",X"A6",X"88",X"4F",X"81",X"02",X"25",X"27",X"AE",X"88",X"1A",X"26",X"F4",X"BE",X"B0",
		X"09",X"27",X"0A",X"A6",X"88",X"4F",X"27",X"18",X"AE",X"88",X"1A",X"26",X"F6",X"BE",X"B0",X"41",
		X"27",X"14",X"A6",X"88",X"4F",X"81",X"02",X"25",X"07",X"AE",X"88",X"1A",X"26",X"F4",X"20",X"06",
		X"AF",X"C8",X"4E",X"6C",X"88",X"4F",X"39",X"8E",X"2E",X"05",X"AF",X"C8",X"3E",X"A6",X"C8",X"30",
		X"E6",X"C8",X"32",X"BD",X"67",X"5E",X"A7",X"C8",X"38",X"27",X"08",X"A7",X"C8",X"16",X"8E",X"2D",
		X"06",X"AF",X"4A",X"7E",X"2F",X"69",X"A6",X"C8",X"16",X"8E",X"2F",X"B2",X"AE",X"86",X"A6",X"C8",
		X"30",X"E6",X"C8",X"32",X"6E",X"84",X"10",X"A3",X"C8",X"5E",X"27",X"08",X"20",X"12",X"10",X"A3",
		X"C8",X"5E",X"26",X"14",X"BD",X"F9",X"16",X"39",X"C1",X"EC",X"25",X"5D",X"C6",X"EC",X"20",X"3F",
		X"C1",X"B1",X"22",X"55",X"C6",X"B1",X"20",X"27",X"C1",X"38",X"25",X"04",X"C6",X"38",X"20",X"2F",
		X"C1",X"36",X"22",X"45",X"C6",X"36",X"20",X"17",X"C1",X"35",X"22",X"3D",X"C6",X"35",X"20",X"0F",
		X"C1",X"97",X"22",X"35",X"C6",X"98",X"8E",X"00",X"00",X"AF",X"C8",X"34",X"BD",X"39",X"2F",X"E7",
		X"C8",X"32",X"EC",X"C8",X"36",X"2A",X"22",X"CC",X"00",X"00",X"ED",X"C8",X"36",X"20",X"1A",X"E7",
		X"C8",X"32",X"EC",X"C8",X"36",X"2F",X"12",X"20",X"EE",X"C1",X"68",X"25",X"0C",X"C6",X"68",X"20",
		X"EE",X"C1",X"48",X"25",X"04",X"C6",X"48",X"20",X"E6",X"CC",X"2C",X"0C",X"ED",X"4A",X"39",X"A7",
		X"C8",X"30",X"EC",X"C8",X"34",X"2A",X"F2",X"CC",X"00",X"00",X"ED",X"C8",X"34",X"20",X"EA",X"A7",
		X"C8",X"30",X"EC",X"C8",X"34",X"2F",X"E2",X"20",X"EE",X"81",X"24",X"22",X"DC",X"86",X"24",X"20",
		X"DE",X"81",X"70",X"25",X"D4",X"86",X"70",X"20",X"E6",X"81",X"1E",X"22",X"CC",X"86",X"1E",X"20",
		X"CE",X"81",X"73",X"25",X"C4",X"86",X"73",X"20",X"D6",X"81",X"27",X"22",X"BC",X"86",X"27",X"20",
		X"BE",X"81",X"6C",X"25",X"B4",X"86",X"6C",X"20",X"C6",X"81",X"29",X"22",X"AC",X"86",X"29",X"20",
		X"AE",X"81",X"6A",X"25",X"A4",X"86",X"6A",X"20",X"B6",X"C6",X"10",X"E7",X"C8",X"14",X"E6",X"C8",
		X"32",X"E7",X"C8",X"15",X"86",X"01",X"20",X"97",X"C6",X"80",X"E7",X"C8",X"14",X"E6",X"C8",X"32",
		X"E7",X"C8",X"15",X"20",X"9A",X"8E",X"2E",X"80",X"AF",X"C8",X"3E",X"A6",X"C8",X"48",X"BB",X"A8",
		X"F9",X"A7",X"C8",X"48",X"24",X"0B",X"6C",X"C8",X"47",X"6A",X"C8",X"3C",X"2A",X"03",X"6F",X"C8",
		X"3C",X"EC",X"C8",X"36",X"2D",X"23",X"26",X"17",X"EC",X"C8",X"34",X"26",X"2A",X"6C",X"C8",X"4A",
		X"A6",X"C8",X"4A",X"81",X"08",X"25",X"46",X"BD",X"39",X"2F",X"6F",X"C8",X"4A",X"20",X"3E",X"E3",
		X"C8",X"32",X"A1",X"C8",X"5F",X"22",X"0A",X"20",X"0B",X"E3",X"C8",X"32",X"A1",X"C8",X"5F",X"24",
		X"03",X"A6",X"C8",X"5F",X"ED",X"C8",X"32",X"6F",X"C8",X"4A",X"EC",X"C8",X"34",X"2D",X"0C",X"27",
		X"1C",X"E3",X"C8",X"30",X"A1",X"C8",X"5E",X"22",X"0E",X"20",X"0F",X"E3",X"C8",X"30",X"A1",X"C8",
		X"5E",X"25",X"04",X"81",X"F0",X"25",X"03",X"A6",X"C8",X"5E",X"ED",X"C8",X"30",X"7E",X"2F",X"69",
		X"8E",X"2F",X"5B",X"AF",X"C8",X"3E",X"EC",X"C8",X"34",X"2D",X"5F",X"2E",X"30",X"A6",X"C8",X"42",
		X"27",X"18",X"2E",X"04",X"86",X"02",X"20",X"01",X"4F",X"A7",X"C8",X"45",X"6F",X"C8",X"42",X"86",
		X"FF",X"A7",X"C8",X"44",X"CC",X"2F",X"6A",X"7E",X"2F",X"18",X"A6",X"C8",X"45",X"8B",X"FE",X"2A",
		X"02",X"86",X"02",X"A7",X"C8",X"45",X"8E",X"2F",X"76",X"EC",X"86",X"20",X"58",X"A6",X"C8",X"44",
		X"27",X"0F",X"6F",X"C8",X"44",X"86",X"01",X"A7",X"C8",X"42",X"86",X"06",X"A7",X"C8",X"45",X"20",
		X"47",X"A6",X"C8",X"45",X"8B",X"FE",X"2A",X"08",X"8E",X"70",X"C9",X"BD",X"6F",X"D3",X"86",X"06",
		X"A7",X"C8",X"45",X"8E",X"2F",X"7A",X"EC",X"86",X"20",X"2B",X"A6",X"C8",X"44",X"27",X"0F",X"6F",
		X"C8",X"44",X"86",X"FF",X"A7",X"C8",X"42",X"86",X"06",X"A7",X"C8",X"45",X"20",X"1A",X"A6",X"C8",
		X"45",X"8B",X"FE",X"2A",X"08",X"8E",X"70",X"C9",X"BD",X"6F",X"D3",X"86",X"06",X"A7",X"C8",X"45",
		X"8E",X"2F",X"94",X"EC",X"86",X"ED",X"C8",X"40",X"A6",X"C8",X"32",X"81",X"A0",X"22",X"08",X"81",
		X"58",X"22",X"07",X"86",X"04",X"20",X"05",X"4F",X"20",X"02",X"86",X"02",X"AE",X"C8",X"40",X"AE",
		X"86",X"AF",X"42",X"8E",X"2F",X"AE",X"AE",X"86",X"AF",X"46",X"A6",X"46",X"44",X"40",X"AB",X"C8",
		X"30",X"A7",X"44",X"86",X"2A",X"E6",X"C8",X"31",X"2D",X"02",X"86",X"0A",X"A7",X"40",X"A6",X"47",
		X"44",X"40",X"AB",X"C8",X"32",X"A7",X"45",X"6C",X"4F",X"20",X"0E",X"6A",X"C8",X"3B",X"2A",X"09",
		X"A6",X"C8",X"3C",X"A7",X"C8",X"3B",X"7E",X"2C",X"0F",X"39",X"46",X"45",X"4E",X"01",X"53",X"7D",
		X"4A",X"23",X"50",X"BF",X"55",X"4B",X"2F",X"70",X"2F",X"6A",X"2F",X"82",X"2F",X"8E",X"2F",X"82",
		X"2F",X"88",X"46",X"45",X"4E",X"01",X"53",X"7D",X"47",X"8F",X"4E",X"EB",X"54",X"17",X"48",X"D9",
		X"4F",X"D5",X"54",X"B1",X"2F",X"9C",X"2F",X"A8",X"2F",X"9C",X"2F",X"A2",X"4A",X"23",X"50",X"BF",
		X"55",X"4B",X"4B",X"6D",X"51",X"A9",X"55",X"E5",X"4C",X"B7",X"52",X"93",X"56",X"7F",X"0B",X"1E",
		X"09",X"1A",X"07",X"16",X"2D",X"38",X"2D",X"40",X"2D",X"48",X"2D",X"40",X"2D",X"38",X"2D",X"30",
		X"2D",X"30",X"2D",X"48",X"2D",X"48",X"2D",X"16",X"2D",X"16",X"2D",X"C9",X"2D",X"D1",X"2D",X"1E",
		X"2D",X"1E",X"2D",X"D9",X"2D",X"E1",X"2D",X"28",X"2D",X"B9",X"2D",X"C1",X"2D",X"38",X"2D",X"48",
		X"2D",X"40",X"2D",X"A9",X"2D",X"B1",X"2D",X"30",X"2D",X"50",X"2D",X"79",X"2D",X"81",X"2D",X"E9",
		X"2D",X"F8",X"EE",X"E4",X"37",X"36",X"EF",X"E4",X"B7",X"A6",X"06",X"F7",X"A6",X"0A",X"31",X"A5",
		X"10",X"BF",X"A6",X"0B",X"10",X"8E",X"A6",X"11",X"6F",X"A0",X"5A",X"26",X"FB",X"10",X"BF",X"A6",
		X"0D",X"34",X"02",X"4F",X"E6",X"84",X"AA",X"80",X"E7",X"A0",X"6A",X"E4",X"26",X"F6",X"32",X"61",
		X"4D",X"27",X"51",X"10",X"BF",X"A6",X"08",X"31",X"3F",X"10",X"BF",X"A6",X"0F",X"B6",X"A6",X"06",
		X"1F",X"89",X"48",X"48",X"48",X"B7",X"A6",X"05",X"FB",X"A6",X"0A",X"F7",X"A6",X"07",X"1C",X"FE",
		X"CE",X"A6",X"07",X"37",X"12",X"69",X"82",X"4A",X"26",X"FB",X"1C",X"FE",X"37",X"32",X"E6",X"A2",
		X"E2",X"82",X"E7",X"A4",X"4A",X"26",X"F7",X"24",X"12",X"1C",X"FE",X"CE",X"A6",X"0A",X"37",X"32",
		X"E6",X"A2",X"E9",X"82",X"E7",X"A4",X"4A",X"26",X"F7",X"20",X"04",X"6C",X"9F",X"A6",X"0F",X"7A",
		X"A6",X"05",X"26",X"CA",X"BE",X"A6",X"0D",X"10",X"8E",X"A6",X"11",X"39",X"34",X"12",X"A6",X"4C",
		X"81",X"20",X"26",X"02",X"86",X"12",X"8E",X"30",X"8D",X"AD",X"96",X"35",X"92",X"30",X"A1",X"30",
		X"EF",X"30",X"FE",X"30",X"F5",X"30",X"A2",X"31",X"07",X"31",X"0F",X"31",X"0F",X"30",X"CD",X"31",
		X"18",X"39",X"0C",X"71",X"CC",X"00",X"64",X"8E",X"54",X"D3",X"0D",X"38",X"27",X"06",X"CC",X"00",
		X"32",X"8E",X"55",X"23",X"BD",X"32",X"3D",X"D3",X"06",X"DD",X"06",X"8E",X"E2",X"58",X"BF",X"AE",
		X"4F",X"8E",X"70",X"9D",X"BD",X"6F",X"D3",X"8E",X"32",X"78",X"7E",X"31",X"F3",X"A6",X"C8",X"16",
		X"26",X"06",X"CC",X"00",X"32",X"7E",X"31",X"CE",X"BD",X"F9",X"30",X"6C",X"4F",X"86",X"78",X"A7",
		X"4D",X"8E",X"30",X"E7",X"AF",X"4A",X"39",X"6A",X"4D",X"26",X"FB",X"AD",X"D8",X"22",X"39",X"CC",
		X"00",X"32",X"7E",X"31",X"CE",X"CC",X"00",X"4B",X"BD",X"32",X"29",X"7E",X"31",X"CE",X"CC",X"00",
		X"32",X"BD",X"32",X"29",X"7E",X"31",X"CE",X"A6",X"4E",X"2A",X"04",X"BD",X"28",X"17",X"39",X"86",
		X"FF",X"97",X"40",X"8E",X"31",X"4E",X"20",X"03",X"8E",X"31",X"96",X"BD",X"28",X"CC",X"8E",X"31",
		X"42",X"BD",X"28",X"82",X"8E",X"31",X"30",X"AF",X"4A",X"8E",X"70",X"61",X"BD",X"6F",X"D3",X"39",
		X"AD",X"D8",X"47",X"AD",X"D8",X"57",X"A6",X"C8",X"46",X"AA",X"C8",X"56",X"26",X"03",X"AD",X"D8",
		X"22",X"39",X"0A",X"04",X"88",X"04",X"44",X"04",X"22",X"04",X"11",X"00",X"00",X"00",X"01",X"01",
		X"00",X"06",X"01",X"00",X"00",X"01",X"00",X"FA",X"00",X"02",X"01",X"00",X"05",X"01",X"00",X"00",
		X"01",X"00",X"FB",X"00",X"03",X"01",X"00",X"04",X"01",X"00",X"00",X"01",X"00",X"FC",X"00",X"04",
		X"01",X"00",X"03",X"01",X"00",X"00",X"01",X"00",X"FD",X"00",X"05",X"01",X"00",X"02",X"01",X"00",
		X"00",X"01",X"00",X"FE",X"00",X"06",X"01",X"00",X"01",X"01",X"00",X"00",X"01",X"00",X"FF",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"03",X"00",X"01",X"00",X"00",X"01",X"FD",X"00",
		X"00",X"06",X"01",X"02",X"00",X"01",X"00",X"00",X"01",X"FE",X"00",X"00",X"09",X"01",X"01",X"00",
		X"01",X"00",X"00",X"01",X"FF",X"00",X"00",X"07",X"01",X"00",X"00",X"01",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"8E",X"E2",X"58",X"BF",X"AE",X"4F",X"0C",X"71",
		X"D3",X"06",X"DD",X"06",X"8E",X"70",X"99",X"BD",X"6F",X"D3",X"86",X"05",X"A7",X"C8",X"1F",X"A6",
		X"C8",X"32",X"8E",X"32",X"DD",X"81",X"58",X"23",X"0A",X"8E",X"32",X"B9",X"81",X"A0",X"23",X"03",
		X"8E",X"32",X"95",X"AF",X"C8",X"39",X"6F",X"4D",X"8E",X"31",X"FD",X"AF",X"4A",X"6A",X"4D",X"2E",
		X"27",X"AE",X"C8",X"39",X"A6",X"00",X"2A",X"05",X"AD",X"D8",X"22",X"4F",X"39",X"A7",X"4D",X"A6",
		X"C8",X"30",X"E6",X"C8",X"32",X"A3",X"05",X"ED",X"44",X"EC",X"03",X"ED",X"46",X"EC",X"01",X"ED",
		X"42",X"30",X"07",X"AF",X"C8",X"39",X"6C",X"4F",X"39",X"6D",X"C8",X"4E",X"27",X"0E",X"8E",X"E2",
		X"58",X"BF",X"AE",X"4F",X"C3",X"00",X"64",X"8E",X"54",X"D3",X"20",X"01",X"39",X"34",X"46",X"A6",
		X"C8",X"30",X"E6",X"C8",X"32",X"20",X"02",X"34",X"46",X"BD",X"F8",X"AD",X"AF",X"42",X"83",X"04",
		X"0C",X"ED",X"44",X"86",X"14",X"A7",X"4C",X"CC",X"1A",X"22",X"ED",X"40",X"CC",X"82",X"05",X"A7",
		X"4D",X"E7",X"C8",X"1F",X"8E",X"08",X"05",X"AF",X"46",X"8E",X"32",X"70",X"AF",X"4A",X"35",X"C6",
		X"6A",X"4D",X"26",X"03",X"AD",X"D8",X"22",X"39",X"08",X"39",X"2E",X"0B",X"1E",X"05",X"0F",X"0A",
		X"3A",X"78",X"0B",X"1E",X"05",X"0F",X"0A",X"3B",X"C2",X"0B",X"1E",X"05",X"0F",X"0C",X"3D",X"0C",
		X"0B",X"1E",X"05",X"0F",X"FF",X"04",X"37",X"41",X"0F",X"17",X"07",X"0B",X"04",X"38",X"9A",X"0E",
		X"15",X"07",X"0A",X"08",X"39",X"C0",X"12",X"1B",X"09",X"0D",X"0A",X"3B",X"A6",X"0B",X"0E",X"05",
		X"07",X"0A",X"3C",X"40",X"0B",X"0E",X"05",X"07",X"FF",X"04",X"3C",X"DA",X"09",X"0E",X"04",X"07",
		X"04",X"3D",X"58",X"0A",X"0E",X"05",X"07",X"08",X"3D",X"E4",X"0C",X"13",X"06",X"09",X"0A",X"3E",
		X"C8",X"09",X"0B",X"04",X"05",X"0A",X"3F",X"2B",X"09",X"0B",X"04",X"05",X"FF",X"04",X"40",X"2D",
		X"07",X"0A",X"03",X"05",X"04",X"40",X"73",X"07",X"09",X"03",X"04",X"08",X"40",X"B2",X"08",X"0C",
		X"04",X"06",X"0A",X"41",X"12",X"06",X"08",X"03",X"04",X"0A",X"41",X"42",X"06",X"08",X"03",X"04",
		X"FF",X"34",X"76",X"86",X"80",X"B7",X"C5",X"82",X"CC",X"10",X"00",X"BD",X"33",X"87",X"CE",X"E3",
		X"2E",X"BD",X"D4",X"47",X"AE",X"01",X"BD",X"E6",X"B9",X"35",X"F6",X"4F",X"C6",X"80",X"FD",X"C5",
		X"81",X"20",X"13",X"7F",X"C5",X"82",X"BD",X"33",X"87",X"20",X"0B",X"86",X"80",X"B7",X"C5",X"82",
		X"CC",X"10",X"00",X"BD",X"33",X"87",X"BD",X"E6",X"B9",X"CC",X"01",X"10",X"20",X"19",X"7F",X"C5",
		X"82",X"BD",X"33",X"87",X"20",X"0B",X"86",X"80",X"B7",X"C5",X"82",X"CC",X"10",X"00",X"BD",X"33",
		X"87",X"BD",X"E6",X"AB",X"CC",X"FF",X"F0",X"DD",X"AA",X"B6",X"C5",X"82",X"BB",X"C5",X"81",X"B7",
		X"C5",X"80",X"10",X"8E",X"34",X"46",X"8D",X"2D",X"0D",X"AB",X"2B",X"02",X"8D",X"41",X"C6",X"40",
		X"D7",X"A9",X"D7",X"DC",X"BD",X"E5",X"1F",X"B6",X"C5",X"80",X"BD",X"33",X"FE",X"0A",X"A9",X"2A",
		X"F3",X"BD",X"E5",X"1F",X"0F",X"A9",X"39",X"34",X"16",X"B7",X"C5",X"81",X"58",X"9E",X"86",X"3A",
		X"BF",X"C5",X"83",X"35",X"96",X"CE",X"BC",X"DD",X"8E",X"C1",X"00",X"8D",X"37",X"8E",X"C2",X"20",
		X"8D",X"48",X"33",X"41",X"8E",X"C3",X"40",X"8D",X"2B",X"8E",X"C4",X"60",X"8D",X"3C",X"39",X"34",
		X"01",X"1A",X"50",X"7F",X"CB",X"A0",X"8E",X"BC",X"DD",X"BF",X"C8",X"84",X"B6",X"C5",X"80",X"C6",
		X"02",X"FD",X"C8",X"86",X"CC",X"00",X"10",X"B7",X"C8",X"81",X"F7",X"C8",X"80",X"86",X"01",X"B7",
		X"CB",X"A0",X"35",X"81",X"B6",X"C5",X"80",X"34",X"42",X"E6",X"C1",X"54",X"54",X"54",X"54",X"E6",
		X"A5",X"4F",X"ED",X"81",X"6A",X"E4",X"26",X"F1",X"35",X"C2",X"B6",X"C5",X"80",X"34",X"42",X"E6",
		X"C1",X"C4",X"0F",X"E6",X"A5",X"4F",X"ED",X"81",X"6A",X"E4",X"26",X"F3",X"35",X"C2",X"8E",X"34",
		X"26",X"D6",X"A9",X"C4",X"03",X"58",X"58",X"58",X"3A",X"EE",X"81",X"10",X"AE",X"81",X"E6",X"A4",
		X"EB",X"21",X"E7",X"A1",X"24",X"0A",X"E6",X"C4",X"EB",X"94",X"E7",X"C1",X"4A",X"26",X"EF",X"39",
		X"33",X"42",X"4A",X"26",X"E9",X"39",X"BC",X"DE",X"C3",X"40",X"BF",X"AB",X"00",X"00",X"BC",X"DD",
		X"C2",X"20",X"BF",X"AA",X"00",X"00",X"BC",X"DD",X"C1",X"00",X"BF",X"AB",X"00",X"00",X"BC",X"DE",
		X"C4",X"60",X"BF",X"AA",X"00",X"00",X"00",X"10",X"20",X"30",X"40",X"50",X"60",X"70",X"80",X"90",
		X"A0",X"B0",X"C0",X"D0",X"E0",X"F0",X"0D",X"9A",X"27",X"10",X"0A",X"9A",X"26",X"0C",X"CE",X"90",
		X"00",X"BD",X"34",X"6E",X"CE",X"90",X"60",X"BD",X"34",X"6E",X"39",X"BD",X"F9",X"4B",X"EE",X"C8",
		X"12",X"26",X"F8",X"39",X"34",X"01",X"1A",X"50",X"96",X"39",X"10",X"26",X"00",X"B2",X"DC",X"DD",
		X"C3",X"00",X"01",X"DD",X"DD",X"10",X"A3",X"9F",X"BF",X"DF",X"25",X"20",X"96",X"96",X"26",X"19",
		X"DE",X"DF",X"33",X"42",X"37",X"36",X"DF",X"DF",X"BD",X"63",X"61",X"EC",X"9F",X"BF",X"DF",X"10",
		X"83",X"FF",X"FF",X"10",X"26",X"00",X"89",X"97",X"D3",X"7E",X"35",X"30",X"BD",X"39",X"52",X"27",
		X"11",X"A6",X"4E",X"10",X"26",X"00",X"79",X"A6",X"C8",X"38",X"8E",X"35",X"45",X"AD",X"96",X"7E",
		X"35",X"30",X"BD",X"39",X"24",X"27",X"24",X"A6",X"4E",X"26",X"65",X"A6",X"C8",X"27",X"27",X"0E",
		X"AE",X"C8",X"25",X"AF",X"C8",X"14",X"6F",X"C8",X"1D",X"6F",X"C8",X"27",X"20",X"52",X"96",X"F4",
		X"26",X"4E",X"A6",X"4C",X"8E",X"35",X"33",X"AD",X"96",X"20",X"45",X"96",X"D0",X"27",X"07",X"0A",
		X"D0",X"26",X"03",X"BD",X"3D",X"49",X"DC",X"DD",X"10",X"83",X"15",X"18",X"24",X"16",X"96",X"D3",
		X"27",X"2E",X"96",X"65",X"26",X"14",X"96",X"D4",X"26",X"10",X"A6",X"9F",X"BA",X"9D",X"26",X"0A",
		X"96",X"40",X"26",X"06",X"86",X"FF",X"97",X"38",X"20",X"16",X"96",X"D1",X"26",X"0A",X"96",X"D5",
		X"84",X"7F",X"8B",X"80",X"97",X"D1",X"20",X"08",X"0A",X"D1",X"26",X"04",X"86",X"FF",X"97",X"D2",
		X"35",X"81",X"39",X"37",X"07",X"37",X"07",X"35",X"B7",X"35",X"C0",X"36",X"03",X"36",X"61",X"36",
		X"74",X"36",X"9C",X"36",X"74",X"37",X"CA",X"37",X"72",X"37",X"77",X"37",X"7C",X"37",X"81",X"37",
		X"86",X"37",X"8B",X"37",X"90",X"37",X"95",X"37",X"9A",X"37",X"9F",X"37",X"A4",X"37",X"A9",X"37",
		X"AE",X"37",X"B3",X"37",X"B8",X"37",X"CB",X"37",X"D0",X"37",X"D5",X"37",X"DC",X"37",X"E1",X"37",
		X"E6",X"37",X"FA",X"37",X"FF",X"38",X"10",X"38",X"15",X"38",X"1A",X"38",X"1F",X"37",X"E6",X"37",
		X"E6",X"38",X"30",X"38",X"38",X"34",X"02",X"BE",X"B0",X"41",X"BD",X"63",X"28",X"A6",X"88",X"30",
		X"A1",X"C8",X"30",X"26",X"0D",X"A6",X"88",X"32",X"A1",X"C8",X"32",X"26",X"05",X"86",X"FF",X"A7",
		X"88",X"3D",X"35",X"82",X"D6",X"D5",X"4F",X"C3",X"02",X"1C",X"10",X"93",X"DD",X"10",X"24",X"00",
		X"C3",X"CC",X"48",X"38",X"7E",X"36",X"F0",X"86",X"10",X"E6",X"C8",X"56",X"2A",X"39",X"20",X"07",
		X"86",X"20",X"E6",X"C8",X"56",X"2A",X"30",X"A6",X"C8",X"30",X"E6",X"C8",X"32",X"AE",X"C8",X"54",
		X"10",X"A3",X"88",X"14",X"26",X"06",X"96",X"E3",X"81",X"04",X"27",X"06",X"EC",X"88",X"14",X"7E",
		X"36",X"F0",X"A6",X"4C",X"97",X"D4",X"BD",X"38",X"40",X"BD",X"F9",X"4B",X"AE",X"C8",X"54",X"86",
		X"FF",X"A7",X"88",X"50",X"7E",X"37",X"07",X"D6",X"E4",X"26",X"A9",X"D6",X"EA",X"27",X"06",X"8D",
		X"84",X"20",X"02",X"86",X"00",X"B7",X"AF",X"5E",X"AE",X"C8",X"54",X"10",X"27",X"00",X"F8",X"A6",
		X"88",X"30",X"A1",X"88",X"14",X"25",X"12",X"A0",X"88",X"14",X"8D",X"02",X"20",X"14",X"D6",X"D5",
		X"C4",X"7F",X"CB",X"40",X"3D",X"BB",X"AF",X"5E",X"39",X"A6",X"88",X"14",X"A0",X"88",X"30",X"8D",
		X"ED",X"40",X"AB",X"88",X"14",X"34",X"02",X"A6",X"88",X"32",X"A1",X"88",X"15",X"25",X"0F",X"A0",
		X"88",X"15",X"8D",X"02",X"20",X"11",X"D6",X"D6",X"C4",X"7F",X"CB",X"60",X"3D",X"39",X"A6",X"88",
		X"15",X"A0",X"88",X"32",X"8D",X"F0",X"40",X"AB",X"88",X"15",X"1F",X"89",X"35",X"02",X"7E",X"36",
		X"F0",X"96",X"E4",X"26",X"0F",X"AE",X"C8",X"54",X"10",X"27",X"00",X"9B",X"CC",X"20",X"20",X"BD",
		X"37",X"11",X"20",X"7C",X"DC",X"D5",X"84",X"3F",X"C4",X"3F",X"34",X"04",X"A1",X"E0",X"24",X"02",
		X"1E",X"89",X"34",X"02",X"A6",X"C8",X"30",X"81",X"49",X"35",X"02",X"25",X"01",X"40",X"6D",X"C8",
		X"32",X"2E",X"01",X"50",X"AB",X"C8",X"30",X"EB",X"C8",X"32",X"20",X"54",X"A6",X"C8",X"30",X"81",
		X"49",X"2D",X"1F",X"E6",X"C8",X"32",X"C1",X"5C",X"22",X"0C",X"81",X"75",X"22",X"04",X"C6",X"04",
		X"20",X"2D",X"C6",X"06",X"20",X"29",X"C1",X"84",X"22",X"04",X"C6",X"0A",X"20",X"21",X"C6",X"0E",
		X"20",X"1D",X"E6",X"C8",X"32",X"C1",X"5C",X"22",X"0C",X"81",X"20",X"22",X"04",X"C6",X"00",X"20",
		X"0E",X"C6",X"02",X"20",X"0A",X"C1",X"84",X"22",X"04",X"C6",X"08",X"20",X"02",X"C6",X"0C",X"8E",
		X"37",X"30",X"AE",X"85",X"96",X"D5",X"84",X"03",X"A6",X"86",X"8E",X"37",X"60",X"48",X"EC",X"86",
		X"0D",X"96",X"26",X"13",X"34",X"02",X"A6",X"4C",X"81",X"04",X"35",X"02",X"27",X"0A",X"6F",X"C8",
		X"1D",X"6F",X"C8",X"1E",X"ED",X"C8",X"14",X"39",X"ED",X"C8",X"2C",X"86",X"06",X"A7",X"C8",X"2B",
		X"39",X"34",X"06",X"A6",X"88",X"30",X"A0",X"C8",X"30",X"35",X"02",X"2A",X"01",X"40",X"AB",X"C8",
		X"30",X"E6",X"88",X"32",X"E0",X"C8",X"32",X"35",X"04",X"2A",X"01",X"50",X"EB",X"C8",X"32",X"39",
		X"37",X"40",X"37",X"44",X"37",X"48",X"37",X"4C",X"37",X"50",X"37",X"54",X"37",X"58",X"37",X"5C",
		X"01",X"03",X"04",X"08",X"00",X"03",X"04",X"08",X"00",X"01",X"04",X"07",X"00",X"01",X"03",X"07",
		X"03",X"04",X"06",X"08",X"00",X"01",X"05",X"07",X"06",X"08",X"06",X"08",X"05",X"07",X"05",X"07",
		X"12",X"37",X"28",X"37",X"48",X"38",X"67",X"37",X"7E",X"37",X"13",X"B1",X"7E",X"B1",X"28",X"71",
		X"6C",X"71",X"CC",X"31",X"54",X"20",X"44",X"CC",X"31",X"54",X"20",X"3F",X"CC",X"49",X"54",X"20",
		X"3A",X"CC",X"61",X"54",X"20",X"35",X"CC",X"61",X"54",X"20",X"30",X"CC",X"25",X"C4",X"20",X"2B",
		X"CC",X"6D",X"C4",X"20",X"26",X"CC",X"2D",X"54",X"20",X"21",X"CC",X"59",X"54",X"20",X"1C",X"CC",
		X"09",X"C4",X"20",X"17",X"CC",X"85",X"C4",X"20",X"12",X"CC",X"2D",X"74",X"20",X"0D",X"CC",X"61",
		X"74",X"20",X"08",X"CC",X"09",X"3C",X"20",X"03",X"CC",X"85",X"3C",X"0D",X"96",X"26",X"0B",X"ED",
		X"C8",X"14",X"86",X"FF",X"A7",X"C8",X"1E",X"6F",X"C8",X"1D",X"39",X"CC",X"2D",X"74",X"20",X"EB",
		X"CC",X"61",X"74",X"20",X"E6",X"A6",X"C8",X"30",X"C6",X"E4",X"20",X"DF",X"CC",X"25",X"A4",X"20",
		X"DA",X"CC",X"6D",X"A4",X"20",X"D5",X"A6",X"C8",X"30",X"81",X"49",X"25",X"04",X"86",X"65",X"20",
		X"02",X"86",X"31",X"E6",X"C8",X"32",X"CB",X"20",X"20",X"C1",X"CC",X"49",X"54",X"20",X"BC",X"A6",
		X"C8",X"30",X"81",X"49",X"25",X"04",X"86",X"65",X"20",X"02",X"86",X"31",X"C6",X"54",X"20",X"AB",
		X"CC",X"2D",X"54",X"20",X"A6",X"CC",X"65",X"54",X"20",X"A1",X"CC",X"48",X"8C",X"20",X"9C",X"A6",
		X"C8",X"30",X"81",X"49",X"25",X"04",X"86",X"55",X"20",X"02",X"86",X"39",X"C6",X"8C",X"20",X"8B",
		X"86",X"10",X"E6",X"C8",X"32",X"7E",X"37",X"BB",X"86",X"80",X"E6",X"C8",X"32",X"7E",X"37",X"BB",
		X"AE",X"C8",X"4C",X"27",X"0C",X"CC",X"00",X"00",X"ED",X"88",X"4C",X"A7",X"88",X"4B",X"A7",X"88",
		X"4E",X"39",X"96",X"E4",X"27",X"1E",X"A6",X"C8",X"16",X"81",X"06",X"26",X"17",X"AE",X"C8",X"54",
		X"27",X"0E",X"A6",X"C8",X"56",X"27",X"09",X"CC",X"00",X"00",X"ED",X"88",X"54",X"A7",X"88",X"56",
		X"BD",X"F9",X"4B",X"39",X"96",X"D5",X"84",X"7F",X"8B",X"3C",X"A7",X"C8",X"1C",X"8D",X"C1",X"AE",
		X"C8",X"54",X"A6",X"88",X"56",X"2B",X"23",X"6F",X"C8",X"56",X"A6",X"C8",X"30",X"A1",X"88",X"30",
		X"26",X"18",X"E6",X"C8",X"32",X"E1",X"88",X"32",X"26",X"10",X"A6",X"C8",X"16",X"44",X"BD",X"D0",
		X"5E",X"86",X"FF",X"A7",X"C8",X"57",X"86",X"78",X"97",X"D0",X"8E",X"38",X"B0",X"AF",X"4A",X"39",
		X"6A",X"C8",X"1C",X"26",X"5D",X"96",X"96",X"27",X"06",X"8D",X"85",X"BD",X"F9",X"4B",X"39",X"A6",
		X"C8",X"30",X"E6",X"C8",X"32",X"1F",X"01",X"A6",X"C8",X"57",X"2A",X"1D",X"6F",X"4E",X"10",X"AE",
		X"C8",X"54",X"86",X"FF",X"A7",X"A8",X"56",X"86",X"10",X"A7",X"A8",X"42",X"DC",X"D5",X"84",X"0F",
		X"C4",X"0F",X"C3",X"3A",X"5C",X"1F",X"02",X"20",X"1E",X"10",X"AE",X"C8",X"14",X"A6",X"C8",X"30",
		X"81",X"49",X"25",X"06",X"31",X"A9",X"F4",X"00",X"20",X"04",X"31",X"A9",X"0C",X"00",X"8D",X"07",
		X"86",X"FF",X"A7",X"C8",X"1E",X"20",X"0B",X"E6",X"4C",X"A6",X"C8",X"16",X"A7",X"C8",X"17",X"BD",
		X"63",X"B2",X"39",X"34",X"10",X"BE",X"AE",X"F6",X"8C",X"AE",X"92",X"23",X"05",X"EF",X"83",X"BF",
		X"AE",X"F6",X"35",X"90",X"BE",X"AE",X"F6",X"EE",X"81",X"27",X"03",X"BF",X"AE",X"F6",X"39",X"34",
		X"12",X"96",X"39",X"27",X"0E",X"A6",X"4C",X"81",X"04",X"27",X"15",X"81",X"06",X"27",X"11",X"81",
		X"10",X"27",X"0D",X"BE",X"AF",X"5C",X"8C",X"AE",X"F8",X"23",X"05",X"EF",X"83",X"BF",X"AF",X"5C",
		X"35",X"92",X"BE",X"AF",X"5C",X"EE",X"81",X"27",X"03",X"BF",X"AF",X"5C",X"39",X"CC",X"00",X"00",
		X"FD",X"AE",X"F4",X"FD",X"AF",X"5A",X"CE",X"AE",X"F4",X"FF",X"AE",X"F6",X"CE",X"AF",X"5A",X"FF",
		X"AF",X"5C",X"39",X"86",X"01",X"BD",X"E0",X"76",X"8E",X"3C",X"16",X"BD",X"F5",X"42",X"8E",X"3C",
		X"1C",X"BD",X"F5",X"42",X"CC",X"00",X"D2",X"FD",X"AF",X"5F",X"BD",X"E5",X"1F",X"96",X"41",X"85",
		X"04",X"26",X"0D",X"FC",X"AF",X"5F",X"83",X"00",X"01",X"FD",X"AF",X"5F",X"26",X"EC",X"20",X"09",
		X"8E",X"70",X"51",X"BD",X"6F",X"D3",X"BD",X"00",X"82",X"BD",X"E0",X"EC",X"39",X"CE",X"3B",X"99",
		X"10",X"8E",X"AF",X"61",X"8E",X"00",X"0D",X"BD",X"7F",X"33",X"DC",X"10",X"BD",X"65",X"F9",X"8E",
		X"AF",X"69",X"BD",X"66",X"1A",X"86",X"3A",X"A7",X"80",X"8E",X"3B",X"93",X"BD",X"F5",X"CC",X"BD",
		X"3B",X"0F",X"BD",X"53",X"FB",X"D6",X"E3",X"8E",X"3B",X"A6",X"96",X"E1",X"81",X"01",X"23",X"0E",
		X"81",X"02",X"27",X"05",X"8E",X"3B",X"E2",X"20",X"03",X"8E",X"3B",X"CC",X"C0",X"08",X"58",X"AE",
		X"85",X"BD",X"F5",X"A7",X"96",X"E4",X"27",X"32",X"BD",X"3B",X"0F",X"86",X"14",X"BD",X"E5",X"1F",
		X"4A",X"26",X"FA",X"96",X"E1",X"81",X"02",X"24",X"21",X"81",X"01",X"27",X"0E",X"8E",X"62",X"0A",
		X"BD",X"F5",X"A7",X"BD",X"3B",X"0F",X"8E",X"62",X"23",X"20",X"0C",X"8E",X"62",X"10",X"BD",X"F5",
		X"A7",X"BD",X"3B",X"0F",X"8E",X"62",X"29",X"BD",X"F5",X"A7",X"CC",X"00",X"3C",X"BD",X"3A",X"ED",
		X"39",X"BD",X"3A",X"BB",X"27",X"0D",X"8E",X"65",X"4B",X"BD",X"3B",X"0C",X"8E",X"3C",X"E6",X"BD",
		X"3B",X"07",X"39",X"96",X"00",X"27",X"10",X"96",X"40",X"81",X"FF",X"26",X"05",X"8E",X"3C",X"8E",
		X"20",X"1B",X"8E",X"3C",X"69",X"20",X"16",X"8E",X"64",X"9A",X"B6",X"BB",X"B9",X"27",X"0A",X"8E",
		X"64",X"CF",X"96",X"09",X"27",X"03",X"8E",X"65",X"0D",X"BD",X"3B",X"0C",X"39",X"BD",X"3B",X"07",
		X"39",X"BD",X"3A",X"BB",X"27",X"38",X"8E",X"65",X"79",X"BD",X"3B",X"0C",X"8E",X"3C",X"EC",X"BD",
		X"3B",X"07",X"96",X"71",X"81",X"14",X"25",X"1F",X"8E",X"65",X"91",X"BD",X"3B",X"0C",X"CC",X"01",
		X"F4",X"34",X"01",X"1A",X"50",X"D3",X"06",X"DD",X"06",X"35",X"01",X"8E",X"E2",X"58",X"BF",X"AE",
		X"4F",X"8E",X"70",X"59",X"BD",X"6F",X"D3",X"CC",X"00",X"3C",X"BD",X"3A",X"ED",X"39",X"8E",X"3B",
		X"FA",X"BD",X"3B",X"07",X"8E",X"3B",X"FA",X"BD",X"3B",X"18",X"39",X"96",X"E4",X"27",X"26",X"CE",
		X"3C",X"F2",X"10",X"8E",X"AF",X"61",X"8E",X"00",X"0C",X"BD",X"7F",X"33",X"D6",X"71",X"4F",X"BD",
		X"65",X"F9",X"8E",X"AF",X"6D",X"BD",X"66",X"1A",X"1F",X"12",X"CE",X"3C",X"FE",X"8E",X"00",X"09",
		X"BD",X"7F",X"33",X"86",X"FF",X"39",X"8E",X"65",X"A2",X"BD",X"F5",X"A7",X"39",X"FD",X"AF",X"5F",
		X"8D",X"1D",X"BD",X"E5",X"1F",X"FC",X"AF",X"5F",X"83",X"00",X"01",X"FD",X"AF",X"5F",X"26",X"F2",
		X"8E",X"3B",X"8D",X"BD",X"F4",X"87",X"39",X"BD",X"F5",X"CC",X"20",X"03",X"BD",X"F5",X"A7",X"BD",
		X"E5",X"1F",X"B6",X"BC",X"2D",X"2A",X"F8",X"39",X"34",X"01",X"1A",X"50",X"BD",X"F8",X"AD",X"CC",
		X"24",X"05",X"A7",X"4C",X"E7",X"C8",X"33",X"6F",X"4E",X"AF",X"C8",X"30",X"CC",X"3B",X"33",X"ED",
		X"4A",X"35",X"81",X"B6",X"BC",X"2D",X"2A",X"2B",X"AE",X"C8",X"30",X"EC",X"02",X"44",X"56",X"1F",
		X"98",X"E6",X"04",X"ED",X"42",X"ED",X"44",X"86",X"00",X"A7",X"C8",X"1F",X"CC",X"42",X"09",X"ED",
		X"46",X"E6",X"05",X"E7",X"C8",X"32",X"86",X"1F",X"ED",X"40",X"86",X"10",X"A7",X"4D",X"8E",X"3B",
		X"64",X"AF",X"4A",X"39",X"6A",X"4D",X"26",X"24",X"8E",X"3B",X"6F",X"86",X"FF",X"20",X"15",X"6A",
		X"4D",X"26",X"19",X"6A",X"C8",X"33",X"26",X"06",X"AD",X"D8",X"22",X"6C",X"4F",X"39",X"8E",X"3B",
		X"64",X"A6",X"C8",X"32",X"AF",X"4A",X"A7",X"41",X"86",X"0E",X"A7",X"4D",X"39",X"00",X"00",X"52",
		X"60",X"47",X"60",X"AF",X"61",X"00",X"6D",X"60",X"44",X"4D",X"69",X"73",X"73",X"69",X"6F",X"6E",
		X"20",X"20",X"20",X"20",X"20",X"FF",X"60",X"2D",X"60",X"3A",X"60",X"65",X"60",X"8B",X"60",X"BB",
		X"60",X"F0",X"61",X"29",X"61",X"70",X"61",X"B8",X"62",X"5E",X"60",X"65",X"62",X"8C",X"62",X"BB",
		X"63",X"08",X"61",X"29",X"63",X"37",X"62",X"43",X"63",X"8A",X"63",X"AC",X"63",X"C9",X"62",X"5E",
		X"60",X"65",X"64",X"0C",X"64",X"24",X"64",X"3A",X"64",X"51",X"64",X"7A",X"62",X"43",X"63",X"8A",
		X"63",X"AC",X"63",X"C9",X"62",X"5E",X"63",X"EA",X"64",X"0C",X"64",X"24",X"64",X"3A",X"64",X"51",
		X"64",X"7A",X"62",X"43",X"63",X"8A",X"63",X"AC",X"63",X"C9",X"3C",X"00",X"00",X"55",X"60",X"BB",
		X"4D",X"69",X"73",X"73",X"69",X"6F",X"6E",X"20",X"41",X"63",X"63",X"6F",X"6D",X"70",X"6C",X"69",
		X"73",X"68",X"65",X"64",X"21",X"FF",X"3C",X"22",X"00",X"2B",X"60",X"66",X"3C",X"46",X"00",X"2E",
		X"75",X"66",X"31",X"20",X"47",X"4F",X"42",X"42",X"4C",X"45",X"20",X"61",X"6E",X"64",X"20",X"31",
		X"20",X"47",X"52",X"45",X"4E",X"41",X"44",X"45",X"20",X"70",X"65",X"72",X"20",X"6D",X"69",X"73",
		X"73",X"69",X"6F",X"6E",X"2E",X"FF",X"50",X"72",X"65",X"76",X"65",X"6E",X"74",X"20",X"6D",X"6F",
		X"6E",X"65",X"79",X"20",X"66",X"72",X"6F",X"6D",X"20",X"6C",X"65",X"61",X"76",X"69",X"6E",X"67",
		X"20",X"73",X"63",X"72",X"65",X"65",X"6E",X"2E",X"FF",X"3C",X"6F",X"00",X"5E",X"60",X"55",X"54",
		X"75",X"72",X"6B",X"65",X"79",X"73",X"20",X"73",X"75",X"63",X"63",X"65",X"65",X"64",X"2C",X"20",
		X"2D",X"5C",X"5C",X"54",X"72",X"79",X"20",X"61",X"67",X"61",X"69",X"6E",X"2E",X"FF",X"3C",X"94",
		X"00",X"5E",X"60",X"55",X"54",X"75",X"72",X"6B",X"65",X"79",X"73",X"20",X"73",X"75",X"63",X"63",
		X"65",X"65",X"64",X"2C",X"20",X"2D",X"5C",X"5C",X"42",X"79",X"73",X"74",X"61",X"6E",X"64",X"65",
		X"72",X"20",X"64",X"61",X"6D",X"61",X"67",X"65",X"2E",X"FF",X"3C",X"C0",X"00",X"67",X"77",X"22",
		X"54",X"65",X"72",X"6D",X"69",X"6E",X"61",X"74",X"6F",X"72",X"20",X"31",X"20",X"75",X"70",X"FF",
		X"3C",X"D6",X"00",X"67",X"77",X"22",X"54",X"65",X"72",X"6D",X"69",X"6E",X"61",X"74",X"6F",X"72",
		X"20",X"32",X"20",X"75",X"70",X"FF",X"AF",X"61",X"00",X"58",X"90",X"22",X"AF",X"61",X"00",X"55",
		X"78",X"22",X"59",X"6F",X"75",X"20",X"72",X"6F",X"61",X"73",X"74",X"65",X"64",X"20",X"20",X"74",
		X"75",X"72",X"6B",X"65",X"79",X"73",X"FF",X"4F",X"E6",X"C8",X"14",X"C1",X"49",X"25",X"02",X"86",
		X"80",X"A7",X"C8",X"42",X"EC",X"C8",X"14",X"6D",X"C8",X"42",X"27",X"05",X"83",X"FF",X"03",X"20",
		X"03",X"83",X"04",X"03",X"ED",X"C8",X"4C",X"C3",X"03",X"07",X"ED",X"C8",X"4E",X"8E",X"C0",X"00",
		X"BD",X"3D",X"FE",X"CC",X"00",X"01",X"ED",X"44",X"86",X"76",X"AA",X"C8",X"42",X"A7",X"D8",X"3B",
		X"6F",X"C8",X"3D",X"8E",X"3D",X"48",X"AF",X"4A",X"39",X"34",X"01",X"1A",X"50",X"FE",X"B0",X"59",
		X"27",X"0D",X"8E",X"3E",X"15",X"AF",X"C8",X"39",X"8E",X"3D",X"61",X"AF",X"4A",X"6F",X"4D",X"35",
		X"81",X"86",X"02",X"A7",X"C8",X"3D",X"8D",X"53",X"26",X"0B",X"6F",X"4E",X"86",X"78",X"A7",X"4D",
		X"8E",X"3D",X"76",X"AF",X"4A",X"39",X"86",X"04",X"A7",X"C8",X"3D",X"A6",X"4E",X"27",X"1C",X"8E",
		X"54",X"AB",X"EC",X"C8",X"14",X"C0",X"0A",X"BD",X"32",X"47",X"DC",X"06",X"C3",X"00",X"C8",X"DD",
		X"06",X"86",X"12",X"BD",X"70",X"08",X"8E",X"3E",X"1A",X"20",X"0B",X"6A",X"4D",X"26",X"11",X"86",
		X"FF",X"A7",X"4E",X"8E",X"3E",X"1E",X"AF",X"C8",X"39",X"8E",X"3D",X"B1",X"AF",X"4A",X"6F",X"4D",
		X"39",X"86",X"06",X"A7",X"C8",X"3D",X"8D",X"03",X"27",X"86",X"39",X"6A",X"4D",X"2E",X"14",X"AE",
		X"C8",X"39",X"EC",X"81",X"2A",X"02",X"4F",X"39",X"A7",X"4D",X"EA",X"C8",X"42",X"E7",X"D8",X"3B",
		X"AF",X"C8",X"39",X"39",X"A6",X"C8",X"3D",X"8E",X"3D",X"DC",X"6E",X"96",X"3D",X"FA",X"3D",X"E4",
		X"3D",X"E4",X"3D",X"EC",X"8E",X"3E",X"1E",X"AF",X"C8",X"39",X"6F",X"4D",X"8E",X"3D",X"F6",X"AF",
		X"4A",X"86",X"FF",X"A7",X"4E",X"39",X"8D",X"C3",X"26",X"03",X"BD",X"F9",X"4B",X"39",X"EC",X"C8",
		X"14",X"54",X"54",X"54",X"54",X"3A",X"C6",X"55",X"3D",X"AB",X"C8",X"14",X"84",X"F0",X"1F",X"89",
		X"3A",X"AF",X"C8",X"3B",X"39",X"0C",X"31",X"01",X"32",X"FF",X"0C",X"33",X"0C",X"32",X"0C",X"31",
		X"01",X"76",X"FF",X"86",X"34",X"8E",X"3E",X"2C",X"BD",X"F9",X"06",X"39",X"8E",X"3E",X"46",X"31",
		X"C8",X"34",X"86",X"0C",X"E6",X"80",X"E7",X"A0",X"4A",X"26",X"F9",X"CC",X"00",X"01",X"ED",X"44",
		X"8E",X"3E",X"52",X"AF",X"4A",X"39",X"0F",X"00",X"6E",X"65",X"C0",X"51",X"07",X"FF",X"EE",X"E5",
		X"C0",X"61",X"30",X"C8",X"34",X"8D",X"06",X"30",X"C8",X"3A",X"8D",X"01",X"39",X"6A",X"00",X"2E",
		X"12",X"86",X"0F",X"A7",X"00",X"EC",X"02",X"63",X"01",X"2B",X"04",X"A7",X"98",X"04",X"39",X"E7",
		X"98",X"04",X"39",X"39",X"BD",X"F9",X"4B",X"39",X"34",X"16",X"B6",X"AF",X"F6",X"4A",X"2A",X"02",
		X"86",X"38",X"B7",X"AF",X"F6",X"48",X"8E",X"AF",X"86",X"EC",X"86",X"DD",X"D5",X"35",X"96",X"34",
		X"36",X"86",X"38",X"8D",X"05",X"4A",X"26",X"FB",X"35",X"B6",X"34",X"02",X"DC",X"D7",X"48",X"58",
		X"8E",X"AF",X"86",X"10",X"AE",X"85",X"34",X"26",X"EC",X"86",X"E3",X"E4",X"DD",X"D5",X"35",X"26",
		X"10",X"9E",X"D5",X"10",X"AF",X"85",X"0A",X"D8",X"2A",X"06",X"C6",X"37",X"D7",X"D8",X"20",X"08",
		X"0A",X"D7",X"2A",X"04",X"86",X"37",X"97",X"D7",X"35",X"82",X"CC",X"18",X"37",X"DD",X"D7",X"8E",
		X"3E",X"EE",X"10",X"8E",X"AF",X"86",X"C6",X"38",X"EE",X"81",X"EF",X"A1",X"5A",X"26",X"F9",X"CC",
		X"00",X"24",X"BD",X"DF",X"C4",X"BD",X"3E",X"8F",X"C3",X"FF",X"FF",X"26",X"F5",X"39",X"00",X"00",
		X"E7",X"00",X"2C",X"00",X"4F",X"00",X"80",X"00",X"04",X"00",X"7A",X"00",X"74",X"00",X"A6",X"00",
		X"40",X"00",X"78",X"00",X"C1",X"00",X"F1",X"00",X"47",X"00",X"65",X"00",X"34",X"00",X"B9",X"00",
		X"D0",X"00",X"4B",X"00",X"D3",X"00",X"E7",X"00",X"C3",X"00",X"89",X"00",X"CE",X"00",X"49",X"00",
		X"31",X"00",X"F5",X"00",X"B1",X"00",X"86",X"FF",X"24",X"FF",X"C0",X"FF",X"98",X"FF",X"EA",X"00",
		X"46",X"FF",X"D6",X"FF",X"E2",X"00",X"84",X"00",X"9E",X"00",X"0E",X"00",X"F2",X"FF",X"94",X"FF",
		X"40",X"FF",X"08",X"FF",X"1A",X"FF",X"0A",X"FF",X"CC",X"FF",X"80",X"FF",X"F0",X"00",X"C4",X"00",
		X"AC",X"FF",X"96",X"FF",X"F2",X"FF",X"50",X"FF",X"3A",X"FF",X"BE",X"FF",X"B8",X"00",X"34",X"01",
		X"1A",X"10",X"86",X"05",X"CE",X"66",X"4B",X"D6",X"E3",X"58",X"33",X"C5",X"10",X"8E",X"B0",X"6C",
		X"8E",X"00",X"02",X"BD",X"DF",X"A0",X"FE",X"B0",X"6C",X"10",X"8E",X"B0",X"6C",X"10",X"9F",X"DF",
		X"8E",X"02",X"C9",X"BD",X"DF",X"A0",X"CE",X"6E",X"D3",X"C6",X"0D",X"0D",X"E4",X"26",X"02",X"D6",
		X"E1",X"58",X"33",X"C5",X"10",X"8E",X"B1",X"FE",X"8E",X"00",X"02",X"BD",X"DF",X"A0",X"FE",X"B1",
		X"FE",X"10",X"8E",X"B1",X"FE",X"8E",X"00",X"3E",X"BD",X"DF",X"A0",X"35",X"81",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"28",X"43",X"29",X"20",X"31",X"39",
		X"38",X"34",X"2C",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",
		X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"FF",X"FF",X"FF",
		X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"28",X"43",X"29",X"20",X"31",X"39",
		X"38",X"34",X"2C",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",
		X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"CC",X"09",X"12",
		X"DD",X"7F",X"CC",X"09",X"12",X"DD",X"81",X"39",X"0F",X"8E",X"DC",X"81",X"D3",X"6D",X"DD",X"7D",
		X"DC",X"6D",X"90",X"7F",X"24",X"01",X"4F",X"D0",X"80",X"24",X"01",X"5F",X"DD",X"7B",X"8E",X"40",
		X"8E",X"AF",X"4A",X"CC",X"2A",X"00",X"ED",X"40",X"86",X"05",X"A7",X"C8",X"1F",X"DC",X"6D",X"E7",
		X"C8",X"32",X"A7",X"C8",X"30",X"83",X"04",X"09",X"ED",X"44",X"CC",X"09",X"14",X"ED",X"46",X"CC",
		X"09",X"25",X"ED",X"C8",X"48",X"CC",X"09",X"D9",X"ED",X"C8",X"4A",X"CC",X"0A",X"8D",X"ED",X"C8",
		X"4C",X"C6",X"04",X"86",X"02",X"ED",X"C8",X"46",X"6F",X"4D",X"BD",X"41",X"10",X"39",X"8E",X"41",
		X"39",X"AF",X"4A",X"BD",X"41",X"10",X"34",X"40",X"BD",X"F8",X"AD",X"CC",X"0A",X"00",X"ED",X"40",
		X"86",X"22",X"A7",X"4C",X"96",X"6E",X"84",X"0F",X"8B",X"F0",X"ED",X"C8",X"32",X"CC",X"48",X"00",
		X"ED",X"C8",X"30",X"E6",X"C8",X"32",X"ED",X"44",X"86",X"05",X"A7",X"C8",X"1F",X"8E",X"42",X"DB",
		X"96",X"6E",X"44",X"44",X"44",X"84",X"FE",X"AE",X"86",X"EC",X"84",X"ED",X"C8",X"36",X"EC",X"02",
		X"ED",X"C8",X"3B",X"EC",X"04",X"A7",X"4D",X"96",X"6D",X"80",X"48",X"34",X"01",X"24",X"01",X"40",
		X"3D",X"44",X"56",X"44",X"56",X"44",X"56",X"44",X"56",X"35",X"01",X"24",X"05",X"43",X"53",X"C3",
		X"00",X"01",X"ED",X"C8",X"34",X"CC",X"42",X"65",X"ED",X"C8",X"40",X"CC",X"42",X"5D",X"ED",X"C8",
		X"39",X"6F",X"C8",X"42",X"6F",X"C8",X"43",X"6F",X"4E",X"CC",X"41",X"C3",X"ED",X"4A",X"35",X"C0",
		X"6A",X"4D",X"2E",X"24",X"A6",X"C8",X"47",X"A7",X"4D",X"A7",X"4F",X"6A",X"C8",X"46",X"2B",X"0E",
		X"27",X"06",X"EC",X"C8",X"48",X"ED",X"42",X"39",X"EC",X"C8",X"4A",X"ED",X"42",X"39",X"EC",X"C8",
		X"4C",X"ED",X"42",X"86",X"02",X"A7",X"C8",X"46",X"39",X"0D",X"8E",X"27",X"09",X"8E",X"41",X"4A",
		X"BD",X"F9",X"33",X"6C",X"4F",X"39",X"BD",X"41",X"10",X"39",X"8E",X"70",X"85",X"BD",X"6F",X"D3",
		X"86",X"05",X"8E",X"41",X"58",X"8D",X"4F",X"39",X"8D",X"22",X"8E",X"41",X"62",X"86",X"09",X"8D",
		X"45",X"39",X"8D",X"2D",X"8E",X"41",X"6C",X"86",X"09",X"8D",X"3B",X"39",X"8D",X"0E",X"8E",X"41",
		X"76",X"86",X"09",X"8D",X"31",X"39",X"8D",X"19",X"AD",X"D8",X"22",X"39",X"8E",X"90",X"00",X"BD",
		X"45",X"45",X"27",X"0C",X"10",X"8E",X"BF",X"7B",X"BD",X"46",X"34",X"26",X"FB",X"BD",X"45",X"56",
		X"39",X"8E",X"90",X"60",X"BD",X"45",X"45",X"27",X"0C",X"10",X"8E",X"BF",X"7B",X"BD",X"46",X"34",
		X"26",X"FB",X"BD",X"45",X"56",X"39",X"A7",X"4D",X"AF",X"C8",X"40",X"8E",X"41",X"B1",X"AF",X"4A",
		X"39",X"6A",X"4D",X"26",X"05",X"AE",X"C8",X"40",X"AF",X"4A",X"39",X"A6",X"4E",X"26",X"03",X"BD",
		X"28",X"1B",X"39",X"6A",X"4D",X"26",X"10",X"03",X"8E",X"6C",X"4E",X"8E",X"42",X"86",X"AF",X"C8",
		X"39",X"8E",X"42",X"53",X"AF",X"4A",X"39",X"6A",X"C8",X"43",X"2E",X"10",X"AE",X"C8",X"40",X"A6",
		X"80",X"A7",X"C8",X"43",X"EC",X"81",X"ED",X"C8",X"44",X"AF",X"C8",X"40",X"6A",X"C8",X"42",X"2E",
		X"27",X"AE",X"C8",X"39",X"EC",X"81",X"26",X"04",X"AE",X"84",X"EC",X"1E",X"AF",X"C8",X"39",X"A7",
		X"C8",X"42",X"AE",X"C8",X"44",X"3A",X"EC",X"81",X"ED",X"42",X"EC",X"84",X"ED",X"46",X"54",X"E7",
		X"C8",X"3F",X"5F",X"44",X"56",X"ED",X"C8",X"3D",X"EC",X"C8",X"37",X"A3",X"C8",X"3B",X"ED",X"C8",
		X"37",X"A6",X"C8",X"36",X"82",X"00",X"A7",X"C8",X"36",X"EC",X"C8",X"32",X"A3",X"C8",X"36",X"ED",
		X"C8",X"32",X"A0",X"C8",X"3F",X"A7",X"45",X"EC",X"C8",X"30",X"E3",X"C8",X"34",X"ED",X"C8",X"30",
		X"A3",X"C8",X"3D",X"A7",X"44",X"A6",X"40",X"84",X"DF",X"5D",X"2A",X"02",X"8A",X"20",X"A7",X"40",
		X"6C",X"4F",X"39",X"BD",X"31",X"FD",X"26",X"04",X"96",X"43",X"97",X"42",X"39",X"0A",X"00",X"0A",
		X"04",X"00",X"00",X"42",X"5F",X"14",X"42",X"6E",X"1E",X"42",X"76",X"78",X"42",X"7E",X"13",X"E1",
		X"05",X"08",X"14",X"09",X"04",X"08",X"14",X"29",X"04",X"07",X"14",X"45",X"04",X"07",X"14",X"61",
		X"03",X"05",X"14",X"70",X"03",X"06",X"02",X"41",X"72",X"13",X"25",X"09",X"12",X"04",X"44",X"31",
		X"13",X"25",X"09",X"12",X"04",X"46",X"F0",X"13",X"25",X"09",X"12",X"04",X"49",X"AF",X"13",X"25",
		X"09",X"12",X"04",X"4C",X"6E",X"13",X"25",X"09",X"12",X"02",X"41",X"72",X"13",X"25",X"09",X"12",
		X"04",X"44",X"31",X"13",X"25",X"09",X"12",X"04",X"46",X"F0",X"13",X"25",X"09",X"12",X"04",X"49",
		X"AF",X"13",X"25",X"09",X"12",X"04",X"4C",X"6E",X"13",X"25",X"09",X"12",X"04",X"4F",X"2D",X"13",
		X"25",X"09",X"12",X"04",X"51",X"EC",X"13",X"25",X"09",X"12",X"FF",X"42",X"FB",X"43",X"01",X"43",
		X"07",X"43",X"0D",X"43",X"13",X"43",X"19",X"43",X"1F",X"43",X"25",X"43",X"2B",X"43",X"31",X"43",
		X"37",X"43",X"3D",X"43",X"43",X"43",X"49",X"43",X"4F",X"43",X"55",X"06",X"E8",X"19",X"13",X"47",
		X"3A",X"08",X"B5",X"27",X"B3",X"47",X"3A",X"08",X"AF",X"29",X"32",X"47",X"3A",X"0A",X"0F",X"37",
		X"22",X"42",X"3F",X"0A",X"A0",X"3D",X"6D",X"42",X"3F",X"0B",X"1C",X"43",X"1B",X"42",X"3F",X"0B",
		X"CC",X"4E",X"E0",X"3D",X"44",X"0C",X"3E",X"54",X"D7",X"3D",X"44",X"0B",X"3E",X"4E",X"B2",X"3D",
		X"44",X"0B",X"A3",X"54",X"42",X"3D",X"44",X"0D",X"9F",X"78",X"A7",X"33",X"51",X"0D",X"37",X"77",
		X"CE",X"33",X"51",X"0B",X"F8",X"6E",X"89",X"33",X"51",X"0A",X"B7",X"65",X"27",X"33",X"51",X"0A",
		X"44",X"63",X"D5",X"33",X"51",X"08",X"24",X"51",X"82",X"33",X"51",X"34",X"01",X"1A",X"50",X"BD",
		X"00",X"CC",X"BD",X"F8",X"AD",X"CC",X"04",X"1E",X"97",X"37",X"E7",X"4C",X"CC",X"50",X"11",X"ED",
		X"40",X"CC",X"01",X"01",X"ED",X"46",X"8E",X"43",X"97",X"AF",X"4A",X"BD",X"44",X"69",X"ED",X"C8",
		X"14",X"E7",X"C8",X"32",X"5F",X"ED",X"C8",X"30",X"0F",X"9E",X"35",X"81",X"BD",X"00",X"D6",X"BD",
		X"F9",X"4B",X"0F",X"42",X"0F",X"39",X"39",X"96",X"9E",X"26",X"FB",X"BD",X"44",X"69",X"ED",X"C8",
		X"14",X"A6",X"C8",X"15",X"A0",X"C8",X"32",X"BD",X"44",X"AF",X"E3",X"C8",X"32",X"ED",X"C8",X"32",
		X"A6",X"C8",X"14",X"5F",X"A3",X"C8",X"30",X"34",X"06",X"2A",X"05",X"43",X"53",X"C3",X"00",X"01",
		X"81",X"0F",X"35",X"06",X"22",X"09",X"58",X"49",X"BD",X"44",X"AF",X"47",X"56",X"47",X"56",X"E3",
		X"C8",X"30",X"81",X"8F",X"23",X"02",X"86",X"8F",X"ED",X"C8",X"30",X"E6",X"C8",X"32",X"DD",X"3B",
		X"ED",X"44",X"CC",X"50",X"F0",X"6D",X"C8",X"31",X"2A",X"03",X"CC",X"90",X"0F",X"A7",X"40",X"D7",
		X"72",X"6C",X"4F",X"96",X"41",X"85",X"01",X"27",X"22",X"D6",X"42",X"26",X"1E",X"8E",X"70",X"89",
		X"BD",X"6F",X"D3",X"03",X"42",X"BD",X"00",X"D6",X"CC",X"EC",X"EB",X"DD",X"1D",X"DC",X"3B",X"DD",
		X"6D",X"8E",X"40",X"38",X"86",X"16",X"BD",X"F8",X"FE",X"96",X"41",X"85",X"02",X"27",X"17",X"D6",
		X"52",X"27",X"13",X"8E",X"70",X"6D",X"BD",X"6F",X"D3",X"0F",X"52",X"D6",X"3F",X"D7",X"39",X"CC",
		X"ED",X"10",X"DD",X"1F",X"96",X"41",X"94",X"37",X"26",X"0B",X"96",X"9B",X"94",X"E4",X"27",X"04",
		X"0A",X"5F",X"27",X"0D",X"39",X"BD",X"00",X"82",X"86",X"1E",X"8E",X"70",X"95",X"0F",X"B4",X"20",
		X"08",X"BD",X"00",X"A2",X"86",X"06",X"8E",X"70",X"8D",X"97",X"5F",X"0F",X"37",X"BD",X"6F",X"D3",
		X"8E",X"44",X"EC",X"86",X"26",X"BD",X"F8",X"FE",X"39",X"96",X"E7",X"27",X"03",X"DC",X"E5",X"39",
		X"8E",X"47",X"0D",X"96",X"4E",X"84",X"3F",X"A6",X"86",X"80",X"00",X"2E",X"01",X"4F",X"C6",X"77",
		X"3D",X"58",X"49",X"58",X"49",X"58",X"49",X"C3",X"10",X"80",X"81",X"F0",X"23",X"02",X"86",X"F0",
		X"34",X"02",X"96",X"4F",X"84",X"3F",X"A6",X"86",X"80",X"04",X"2E",X"01",X"4F",X"C6",X"AD",X"3D",
		X"58",X"49",X"58",X"49",X"C3",X"02",X"80",X"81",X"8F",X"23",X"02",X"86",X"8F",X"35",X"84",X"C6",
		X"00",X"8E",X"44",X"CC",X"24",X"0E",X"40",X"81",X"0F",X"22",X"03",X"48",X"EC",X"86",X"43",X"53",
		X"C3",X"00",X"01",X"39",X"81",X"0F",X"22",X"03",X"48",X"EC",X"86",X"39",X"00",X"00",X"00",X"08",
		X"00",X"10",X"00",X"20",X"00",X"40",X"01",X"00",X"03",X"00",X"04",X"00",X"05",X"00",X"06",X"00",
		X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"96",X"73",X"A7",X"4D",
		X"8E",X"44",X"F6",X"AF",X"4A",X"39",X"6A",X"4D",X"26",X"21",X"86",X"04",X"97",X"37",X"8E",X"90",
		X"00",X"8D",X"42",X"27",X"17",X"8D",X"31",X"10",X"8E",X"BF",X"75",X"BD",X"46",X"3C",X"8D",X"46",
		X"10",X"2E",X"01",X"3E",X"2B",X"1C",X"8E",X"45",X"1C",X"AF",X"4A",X"39",X"8E",X"90",X"60",X"8D",
		X"24",X"27",X"0F",X"8D",X"13",X"10",X"8E",X"BF",X"75",X"BD",X"46",X"3C",X"8D",X"28",X"10",X"2E",
		X"01",X"20",X"8E",X"46",X"BD",X"AF",X"4A",X"39",X"DC",X"79",X"D3",X"3B",X"DD",X"77",X"DC",X"3B",
		X"93",X"79",X"DD",X"75",X"39",X"9F",X"61",X"10",X"AE",X"88",X"12",X"27",X"08",X"CC",X"00",X"00",
		X"ED",X"A8",X"10",X"86",X"FF",X"39",X"34",X"01",X"9E",X"61",X"10",X"AE",X"88",X"12",X"AF",X"A8",
		X"10",X"35",X"81",X"34",X"40",X"E6",X"07",X"C0",X"12",X"58",X"58",X"CE",X"45",X"91",X"33",X"C5",
		X"A6",X"88",X"30",X"E6",X"88",X"32",X"A3",X"C4",X"E1",X"23",X"22",X"13",X"81",X"EA",X"22",X"04",
		X"A1",X"22",X"22",X"0B",X"E3",X"42",X"E1",X"21",X"25",X"05",X"A1",X"20",X"25",X"01",X"4F",X"35",
		X"C0",X"02",X"09",X"04",X"0E",X"00",X"00",X"00",X"00",X"02",X"0A",X"04",X"0D",X"03",X"0A",X"05",
		X"0F",X"01",X"0B",X"03",X"03",X"03",X"0B",X"05",X"0F",X"00",X"00",X"00",X"00",X"03",X"0C",X"06",
		X"12",X"01",X"0D",X"03",X"04",X"03",X"0D",X"06",X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"0F",X"04",X"06",X"EC",X"88",X"4C",X"E1",X"23",X"10",X"22",X"00",X"7D",X"A1",X"22",
		X"10",X"22",X"00",X"77",X"EC",X"88",X"4E",X"E1",X"21",X"25",X"70",X"A1",X"20",X"25",X"6C",X"A6",
		X"0E",X"26",X"68",X"86",X"01",X"A7",X"0E",X"35",X"C0",X"EC",X"04",X"E1",X"23",X"22",X"5C",X"81",
		X"EA",X"22",X"04",X"A1",X"22",X"22",X"54",X"E3",X"06",X"E1",X"21",X"23",X"4E",X"A1",X"20",X"23",
		X"4A",X"A6",X"0E",X"26",X"0B",X"BD",X"45",X"63",X"26",X"41",X"86",X"01",X"A7",X"0E",X"35",X"C0",
		X"4F",X"35",X"C0",X"EC",X"04",X"E1",X"23",X"22",X"32",X"A1",X"22",X"22",X"2E",X"E3",X"06",X"E1",
		X"21",X"23",X"28",X"A1",X"20",X"23",X"24",X"A6",X"0E",X"26",X"06",X"86",X"01",X"A7",X"0E",X"35",
		X"C0",X"4F",X"35",X"C0",X"34",X"40",X"CE",X"47",X"93",X"4F",X"20",X"0D",X"34",X"40",X"CE",X"47",
		X"5D",X"86",X"FF",X"20",X"04",X"A6",X"0C",X"6E",X"D6",X"97",X"90",X"AE",X"88",X"10",X"26",X"F5",
		X"35",X"C0",X"AD",X"D8",X"22",X"39",X"EC",X"04",X"E1",X"23",X"22",X"EF",X"81",X"EA",X"22",X"04",
		X"A1",X"22",X"22",X"E7",X"E3",X"06",X"E1",X"21",X"23",X"E1",X"A1",X"20",X"23",X"DD",X"96",X"90",
		X"27",X"05",X"BD",X"D7",X"BA",X"27",X"D4",X"A6",X"0E",X"26",X"0E",X"86",X"01",X"E6",X"0C",X"C1",
		X"0E",X"22",X"02",X"97",X"9E",X"A7",X"0E",X"35",X"C0",X"86",X"FF",X"35",X"C0",X"EC",X"04",X"E1",
		X"23",X"22",X"B8",X"81",X"EA",X"22",X"04",X"A1",X"22",X"22",X"B0",X"E3",X"06",X"E1",X"21",X"23",
		X"AA",X"A1",X"20",X"23",X"A6",X"A6",X"0E",X"26",X"10",X"BD",X"45",X"63",X"26",X"06",X"86",X"01",
		X"A7",X"0E",X"35",X"C0",X"86",X"FF",X"A7",X"88",X"46",X"86",X"FF",X"35",X"C0",X"CC",X"02",X"2A",
		X"A7",X"C8",X"50",X"E7",X"40",X"DC",X"3B",X"83",X"02",X"04",X"ED",X"44",X"CC",X"05",X"09",X"ED",
		X"46",X"8E",X"46",X"DE",X"AF",X"4A",X"8E",X"47",X"4D",X"AF",X"C8",X"39",X"20",X"12",X"6A",X"C8",
		X"50",X"26",X"06",X"8E",X"70",X"91",X"BD",X"6F",X"D3",X"6A",X"4D",X"2E",X"13",X"AE",X"C8",X"39",
		X"A6",X"80",X"2A",X"03",X"6E",X"D8",X"22",X"A7",X"4D",X"EC",X"81",X"ED",X"42",X"AF",X"C8",X"39",
		X"6C",X"4F",X"39",X"86",X"04",X"97",X"73",X"CC",X"00",X"00",X"DD",X"79",X"39",X"00",X"01",X"03",
		X"02",X"07",X"06",X"04",X"05",X"0F",X"0E",X"0C",X"0D",X"08",X"09",X"0B",X"0A",X"1F",X"1E",X"1C",
		X"1D",X"18",X"19",X"1B",X"1A",X"10",X"11",X"13",X"12",X"17",X"16",X"14",X"15",X"3F",X"3E",X"3C",
		X"3D",X"38",X"39",X"3B",X"3A",X"30",X"31",X"33",X"32",X"37",X"36",X"34",X"35",X"20",X"21",X"23",
		X"22",X"27",X"26",X"24",X"25",X"2F",X"2E",X"2C",X"2D",X"28",X"29",X"2B",X"2A",X"06",X"1B",X"99",
		X"04",X"1B",X"C6",X"04",X"1B",X"F3",X"02",X"1C",X"20",X"02",X"1C",X"4D",X"FF",X"46",X"4B",X"46",
		X"13",X"45",X"E9",X"45",X"E9",X"46",X"8D",X"46",X"56",X"46",X"56",X"46",X"56",X"46",X"56",X"46",
		X"56",X"46",X"4B",X"46",X"4B",X"46",X"56",X"46",X"56",X"46",X"56",X"46",X"4B",X"46",X"56",X"46",
		X"4B",X"46",X"4B",X"46",X"4B",X"46",X"4B",X"46",X"4B",X"45",X"C5",X"46",X"56",X"46",X"13",X"46",
		X"4B",X"46",X"4B",X"46",X"4B",X"46",X"13",X"46",X"13",X"46",X"13",X"46",X"13",X"46",X"4B",X"46",
		X"4B",X"46",X"4B",X"46",X"56",X"46",X"56",X"46",X"4B",X"46",X"4B",X"46",X"56",X"46",X"56",X"46",
		X"56",X"46",X"4B",X"46",X"13",X"46",X"4B",X"46",X"4B",X"46",X"4B",X"46",X"4B",X"46",X"4B",X"45",
		X"C5",X"46",X"56",X"46",X"13",X"46",X"4B",X"46",X"4B",X"CC",X"0A",X"00",X"ED",X"40",X"86",X"05",
		X"A7",X"C8",X"1F",X"CC",X"10",X"0E",X"ED",X"46",X"CC",X"01",X"F8",X"ED",X"C8",X"48",X"CC",X"02",
		X"D8",X"ED",X"C8",X"4A",X"CC",X"03",X"B8",X"ED",X"C8",X"4C",X"ED",X"42",X"CC",X"08",X"08",X"E7",
		X"C8",X"3F",X"5F",X"ED",X"C8",X"3D",X"C6",X"02",X"86",X"02",X"ED",X"C8",X"46",X"6F",X"4D",X"8E",
		X"49",X"E8",X"AF",X"C8",X"42",X"6F",X"C8",X"40",X"6F",X"C8",X"1D",X"6F",X"4E",X"0F",X"5C",X"BD",
		X"48",X"65",X"BD",X"48",X"6E",X"39",X"BD",X"41",X"10",X"AD",X"D8",X"50",X"27",X"03",X"8D",X"4E",
		X"39",X"8D",X"4B",X"EC",X"C8",X"36",X"27",X"0F",X"8E",X"48",X"7E",X"96",X"5B",X"81",X"04",X"26",
		X"03",X"8E",X"49",X"C7",X"AF",X"C8",X"4E",X"8E",X"48",X"40",X"AF",X"4A",X"BD",X"48",X"9D",X"39",
		X"A6",X"C8",X"1D",X"27",X"20",X"A6",X"4E",X"10",X"26",X"00",X"DC",X"BD",X"41",X"10",X"8D",X"1E",
		X"96",X"5C",X"27",X"10",X"8E",X"07",X"38",X"AF",X"C8",X"48",X"0A",X"5C",X"26",X"06",X"8E",X"01",
		X"F8",X"AF",X"C8",X"48",X"39",X"BD",X"49",X"58",X"8E",X"48",X"16",X"AF",X"4A",X"39",X"A6",X"C8",
		X"30",X"E6",X"C8",X"32",X"AD",X"D8",X"4E",X"80",X"08",X"C0",X"08",X"ED",X"44",X"39",X"34",X"06",
		X"A6",X"C8",X"52",X"8B",X"0E",X"A7",X"C8",X"52",X"24",X"11",X"A6",X"C8",X"47",X"4C",X"A7",X"C8",
		X"47",X"81",X"07",X"25",X"06",X"8E",X"49",X"E7",X"AF",X"C8",X"4E",X"35",X"86",X"86",X"FF",X"A7",
		X"C8",X"1D",X"EC",X"C8",X"14",X"81",X"AC",X"24",X"05",X"C1",X"00",X"27",X"01",X"39",X"AD",X"D8",
		X"22",X"39",X"EC",X"C8",X"34",X"8D",X"13",X"25",X"03",X"8D",X"28",X"39",X"A6",X"40",X"84",X"DF",
		X"6D",X"C8",X"30",X"2A",X"02",X"8A",X"20",X"A7",X"40",X"39",X"E3",X"C8",X"30",X"A1",X"C8",X"30",
		X"27",X"02",X"6C",X"4F",X"ED",X"C8",X"30",X"8B",X"20",X"E6",X"C8",X"14",X"CB",X"20",X"34",X"04",
		X"A1",X"E0",X"39",X"6C",X"4F",X"A6",X"C8",X"14",X"A7",X"C8",X"30",X"6F",X"C8",X"31",X"39",X"EC",
		X"C8",X"36",X"2B",X"07",X"8D",X"0C",X"25",X"09",X"8D",X"21",X"39",X"8D",X"05",X"22",X"02",X"8D",
		X"1A",X"39",X"E3",X"C8",X"32",X"A1",X"C8",X"32",X"27",X"02",X"6C",X"4F",X"ED",X"C8",X"32",X"8B",
		X"0A",X"E6",X"C8",X"15",X"CB",X"0A",X"34",X"04",X"A1",X"E0",X"39",X"6C",X"4F",X"A6",X"C8",X"15",
		X"A7",X"C8",X"32",X"6F",X"C8",X"33",X"39",X"8E",X"70",X"65",X"BD",X"6F",X"D3",X"86",X"FE",X"97",
		X"40",X"8E",X"00",X"00",X"96",X"5B",X"81",X"04",X"26",X"08",X"86",X"40",X"A7",X"C8",X"15",X"8E",
		X"00",X"CA",X"AF",X"C8",X"36",X"8E",X"49",X"FA",X"AF",X"C8",X"39",X"8E",X"49",X"51",X"AF",X"4A",
		X"39",X"BD",X"48",X"EF",X"BD",X"31",X"FD",X"39",X"EC",X"C8",X"14",X"A1",X"C8",X"30",X"27",X"19",
		X"8E",X"00",X"40",X"AF",X"C8",X"34",X"8E",X"00",X"00",X"AF",X"C8",X"36",X"8E",X"48",X"B2",X"AF",
		X"C8",X"50",X"8E",X"49",X"C7",X"AF",X"C8",X"4E",X"39",X"8E",X"00",X"30",X"E1",X"C8",X"32",X"27",
		X"1B",X"22",X"03",X"8E",X"FF",X"D0",X"AF",X"C8",X"36",X"8E",X"00",X"00",X"AF",X"C8",X"34",X"8E",
		X"48",X"EF",X"AF",X"C8",X"50",X"8E",X"49",X"E7",X"AF",X"C8",X"4E",X"39",X"39",X"A6",X"4E",X"26",
		X"25",X"86",X"02",X"A7",X"C8",X"47",X"EC",X"C8",X"34",X"27",X"0D",X"86",X"AC",X"A7",X"C8",X"14",
		X"8E",X"00",X"C0",X"AF",X"C8",X"34",X"20",X"0B",X"86",X"00",X"A7",X"C8",X"15",X"8E",X"FF",X"A0",
		X"AF",X"C8",X"36",X"6F",X"C8",X"1D",X"39",X"6A",X"C8",X"40",X"2A",X"18",X"6C",X"4F",X"AE",X"C8",
		X"42",X"34",X"06",X"EC",X"81",X"26",X"05",X"8E",X"49",X"E8",X"EC",X"81",X"ED",X"C8",X"40",X"AF",
		X"C8",X"42",X"35",X"06",X"EB",X"C8",X"41",X"39",X"08",X"00",X"08",X"01",X"08",X"02",X"08",X"01",
		X"08",X"00",X"08",X"FF",X"08",X"FE",X"08",X"FF",X"00",X"00",X"14",X"07",X"38",X"10",X"0E",X"08",
		X"08",X"08",X"04",X"98",X"10",X"0E",X"08",X"08",X"08",X"05",X"78",X"10",X"0E",X"08",X"08",X"08",
		X"06",X"58",X"10",X"0E",X"08",X"08",X"FF",X"5F",X"BD",X"E5",X"61",X"BD",X"F0",X"6B",X"BD",X"E0",
		X"EC",X"4F",X"BD",X"66",X"BC",X"CC",X"03",X"84",X"DD",X"55",X"8E",X"E2",X"C4",X"BF",X"AE",X"55",
		X"7F",X"AE",X"57",X"8E",X"4C",X"C6",X"BD",X"13",X"22",X"8E",X"4C",X"7F",X"BD",X"F5",X"42",X"8E",
		X"4C",X"98",X"BD",X"F5",X"42",X"CC",X"02",X"44",X"10",X"8E",X"4C",X"EB",X"BD",X"4A",X"CE",X"CC",
		X"01",X"55",X"10",X"8E",X"4C",X"F2",X"BD",X"4A",X"D6",X"CC",X"01",X"22",X"10",X"8E",X"4C",X"E4",
		X"8D",X"6C",X"96",X"97",X"27",X"22",X"CC",X"22",X"BB",X"FD",X"A6",X"4D",X"BD",X"4B",X"B2",X"BD",
		X"4A",X"C3",X"10",X"8E",X"4C",X"EB",X"CC",X"44",X"CC",X"FD",X"A6",X"4D",X"BD",X"4B",X"C3",X"BD",
		X"DA",X"A3",X"0F",X"97",X"0F",X"9F",X"20",X"1D",X"10",X"8E",X"4C",X"E4",X"96",X"25",X"BD",X"4B",
		X"04",X"B6",X"BB",X"DE",X"BD",X"4B",X"04",X"96",X"26",X"BD",X"4B",X"0F",X"B6",X"BB",X"DF",X"BD",
		X"4B",X"0F",X"BD",X"4A",X"C3",X"BD",X"70",X"28",X"1C",X"AF",X"BD",X"E5",X"1F",X"DC",X"55",X"C3",
		X"FF",X"FF",X"DD",X"55",X"2E",X"F4",X"8E",X"4C",X"D0",X"BD",X"13",X"22",X"8E",X"4C",X"DA",X"BD",
		X"13",X"22",X"39",X"86",X"03",X"BD",X"E0",X"76",X"C6",X"06",X"BD",X"E5",X"61",X"39",X"8D",X"06",
		X"4C",X"A1",X"26",X"23",X"F9",X"39",X"34",X"46",X"F7",X"A6",X"36",X"AD",X"B8",X"02",X"F7",X"A6",
		X"35",X"BF",X"A6",X"33",X"A6",X"E4",X"4A",X"C6",X"06",X"3D",X"EE",X"24",X"33",X"CB",X"E6",X"E4",
		X"4F",X"BD",X"65",X"FE",X"8E",X"A6",X"37",X"BF",X"A6",X"31",X"BD",X"4B",X"26",X"8E",X"A6",X"31",
		X"AD",X"B4",X"35",X"C6",X"27",X"08",X"40",X"8B",X"0B",X"C6",X"BB",X"BD",X"4A",X"D6",X"39",X"27",
		X"14",X"10",X"8E",X"4C",X"EB",X"40",X"8B",X"26",X"81",X"01",X"26",X"04",X"10",X"8E",X"4C",X"F2",
		X"C6",X"CC",X"BD",X"4A",X"D6",X"39",X"34",X"10",X"8D",X"24",X"CC",X"29",X"20",X"ED",X"81",X"37",
		X"06",X"ED",X"81",X"37",X"02",X"C6",X"20",X"ED",X"81",X"E7",X"80",X"37",X"02",X"8D",X"0F",X"37",
		X"02",X"8D",X"0E",X"37",X"02",X"8D",X"0A",X"CC",X"30",X"FF",X"ED",X"81",X"35",X"90",X"7F",X"A6",
		X"4B",X"34",X"02",X"44",X"44",X"44",X"44",X"8D",X"07",X"35",X"02",X"84",X"0F",X"8D",X"01",X"39",
		X"8A",X"30",X"81",X"30",X"26",X"09",X"F6",X"A6",X"4B",X"26",X"04",X"86",X"20",X"20",X"03",X"7C",
		X"A6",X"4B",X"A7",X"80",X"39",X"CE",X"4B",X"90",X"5F",X"81",X"0E",X"59",X"81",X"1A",X"59",X"58",
		X"33",X"C5",X"E6",X"41",X"8E",X"00",X"1C",X"3A",X"A0",X"C4",X"C6",X"08",X"3D",X"CB",X"85",X"39",
		X"1A",X"AC",X"0E",X"56",X"00",X"00",X"02",X"00",X"81",X"05",X"2E",X"05",X"8E",X"00",X"26",X"20",
		X"05",X"8E",X"00",X"9E",X"80",X"05",X"C6",X"0A",X"3D",X"CB",X"28",X"39",X"C6",X"79",X"8E",X"00",
		X"17",X"39",X"CC",X"00",X"00",X"FD",X"A6",X"4F",X"8D",X"1A",X"BD",X"7E",X"73",X"8D",X"15",X"BD",
		X"7E",X"73",X"39",X"CC",X"01",X"08",X"FD",X"A6",X"4F",X"8D",X"10",X"BD",X"7E",X"73",X"8D",X"0B",
		X"BD",X"7E",X"73",X"39",X"CE",X"AA",X"5A",X"96",X"25",X"20",X"05",X"CE",X"AA",X"1D",X"96",X"26",
		X"27",X"29",X"8D",X"2F",X"34",X"06",X"F6",X"A6",X"50",X"27",X"0E",X"86",X"0E",X"7D",X"A6",X"4C",
		X"26",X"02",X"86",X"0F",X"BD",X"70",X"08",X"8D",X"13",X"35",X"06",X"8D",X"3E",X"2A",X"E5",X"7D",
		X"A6",X"50",X"27",X"07",X"BD",X"00",X"B5",X"C6",X"78",X"8D",X"01",X"39",X"BD",X"E5",X"1F",X"5A",
		X"26",X"FA",X"39",X"4A",X"B7",X"A6",X"4C",X"A6",X"26",X"5F",X"BD",X"4A",X"D6",X"34",X"22",X"10",
		X"9E",X"23",X"E6",X"A4",X"E7",X"C4",X"AE",X"21",X"AF",X"41",X"D6",X"03",X"E7",X"43",X"9E",X"04",
		X"AF",X"44",X"35",X"22",X"F6",X"A6",X"4E",X"BD",X"4A",X"D6",X"39",X"7A",X"A6",X"4C",X"2B",X"3E",
		X"5F",X"BD",X"4A",X"D6",X"4A",X"B1",X"A6",X"4F",X"26",X"04",X"10",X"8E",X"4C",X"F2",X"BD",X"4A",
		X"D6",X"C6",X"06",X"34",X"06",X"30",X"5A",X"A6",X"C4",X"E6",X"84",X"A7",X"80",X"E7",X"C0",X"6A",
		X"61",X"26",X"F4",X"33",X"1A",X"35",X"06",X"F6",X"A6",X"4E",X"BD",X"4A",X"D6",X"B1",X"A6",X"4F",
		X"26",X"04",X"10",X"8E",X"4C",X"EB",X"4C",X"F6",X"A6",X"4D",X"BD",X"4A",X"D6",X"4A",X"39",X"4C",
		X"85",X"00",X"5C",X"25",X"11",X"48",X"45",X"52",X"4F",X"45",X"53",X"20",X"46",X"4F",X"52",X"20",
		X"54",X"48",X"45",X"20",X"44",X"41",X"59",X"FF",X"4C",X"9E",X"00",X"1D",X"6C",X"33",X"43",X"48",
		X"49",X"45",X"46",X"20",X"4C",X"55",X"44",X"5A",X"49",X"41",X"27",X"53",X"20",X"45",X"4C",X"49",
		X"54",X"45",X"20",X"54",X"55",X"52",X"4B",X"45",X"59",X"20",X"54",X"45",X"52",X"4D",X"49",X"4E",
		X"41",X"54",X"4F",X"52",X"53",X"FF",X"00",X"08",X"10",X"2E",X"45",X"02",X"05",X"03",X"4C",X"F9",
		X"00",X"08",X"10",X"27",X"45",X"02",X"06",X"14",X"4C",X"F9",X"00",X"08",X"10",X"27",X"45",X"02",
		X"06",X"14",X"4D",X"12",X"F5",X"42",X"4B",X"98",X"AA",X"24",X"0A",X"F5",X"4F",X"4B",X"75",X"A9",
		X"45",X"25",X"F5",X"42",X"4B",X"AC",X"A9",X"45",X"25",X"4D",X"03",X"4D",X"08",X"4D",X"0D",X"00",
		X"00",X"4C",X"F9",X"77",X"88",X"00",X"4D",X"03",X"77",X"99",X"00",X"4D",X"08",X"88",X"99",X"00",
		X"4D",X"0D",X"4D",X"18",X"00",X"00",X"4D",X"12",X"FF",X"FF",X"FF",X"FF",X"00",X"4D",X"18",X"8E",
		X"4E",X"5B",X"E6",X"C8",X"15",X"2B",X"03",X"8E",X"4E",X"3A",X"8D",X"4F",X"BD",X"28",X"48",X"39",
		X"8E",X"4E",X"CD",X"E6",X"C8",X"30",X"2B",X"03",X"8E",X"4E",X"E3",X"8D",X"3E",X"BD",X"28",X"48",
		X"39",X"8E",X"4E",X"94",X"E6",X"C8",X"15",X"C1",X"A0",X"24",X"0A",X"8E",X"4E",X"88",X"C1",X"58",
		X"24",X"03",X"8E",X"4E",X"7C",X"8D",X"24",X"CC",X"00",X"00",X"ED",X"C8",X"3E",X"96",X"EA",X"27",
		X"16",X"BE",X"B0",X"41",X"27",X"11",X"BD",X"63",X"28",X"A6",X"88",X"30",X"A1",X"C8",X"30",X"26",
		X"06",X"AF",X"C8",X"3E",X"EF",X"88",X"3E",X"BD",X"28",X"48",X"39",X"86",X"05",X"A7",X"C8",X"1F",
		X"EC",X"00",X"ED",X"46",X"EC",X"06",X"ED",X"42",X"EC",X"C8",X"14",X"A7",X"C8",X"30",X"E7",X"C8",
		X"32",X"A3",X"02",X"ED",X"44",X"EC",X"04",X"ED",X"C8",X"39",X"EC",X"08",X"ED",X"C8",X"40",X"EC",
		X"0A",X"A7",X"C8",X"46",X"E7",X"C8",X"2A",X"6F",X"4D",X"6F",X"4E",X"8E",X"4D",X"B1",X"AF",X"4A",
		X"39",X"A6",X"4E",X"27",X"12",X"A6",X"C8",X"46",X"BD",X"70",X"08",X"CC",X"00",X"05",X"D3",X"06",
		X"DD",X"06",X"AE",X"C8",X"40",X"AF",X"4A",X"39",X"6A",X"4D",X"2E",X"16",X"AE",X"C8",X"39",X"A6",
		X"84",X"26",X"02",X"AE",X"01",X"A6",X"80",X"A7",X"4D",X"EC",X"81",X"ED",X"42",X"AF",X"C8",X"39",
		X"6C",X"4F",X"39",X"6A",X"4D",X"2E",X"1A",X"AE",X"C8",X"39",X"A6",X"84",X"26",X"06",X"8E",X"4E",
		X"01",X"AF",X"4A",X"39",X"A6",X"80",X"A7",X"4D",X"EC",X"81",X"ED",X"42",X"AF",X"C8",X"39",X"6C",
		X"4F",X"39",X"BD",X"31",X"FD",X"26",X"20",X"AE",X"C8",X"3E",X"27",X"1B",X"63",X"88",X"41",X"EC",
		X"C8",X"14",X"C0",X"06",X"8E",X"55",X"23",X"BD",X"32",X"47",X"CC",X"00",X"32",X"34",X"01",X"1A",
		X"50",X"D3",X"06",X"DD",X"06",X"35",X"01",X"39",X"BD",X"F9",X"4B",X"6C",X"4F",X"39",X"BD",X"F9",
		X"4B",X"6C",X"4F",X"39",X"BD",X"F9",X"4B",X"6C",X"4F",X"39",X"05",X"05",X"03",X"05",X"4E",X"46",
		X"16",X"12",X"4D",X"C8",X"56",X"00",X"05",X"16",X"2B",X"05",X"16",X"44",X"05",X"16",X"5D",X"05",
		X"16",X"44",X"05",X"16",X"2B",X"05",X"16",X"44",X"00",X"4E",X"4C",X"0A",X"0A",X"07",X"0A",X"4E",
		X"67",X"14",X"82",X"4D",X"C8",X"56",X"00",X"05",X"14",X"E6",X"05",X"15",X"4A",X"05",X"15",X"AE",
		X"05",X"15",X"4A",X"05",X"14",X"E6",X"05",X"15",X"4A",X"00",X"4E",X"6D",X"03",X"0C",X"01",X"0C",
		X"4E",X"A0",X"1F",X"19",X"4E",X"02",X"57",X"07",X"04",X"11",X"02",X"11",X"4E",X"AF",X"32",X"60",
		X"4E",X"02",X"57",X"05",X"05",X"13",X"02",X"13",X"4E",X"BE",X"1D",X"64",X"4E",X"02",X"57",X"07",
		X"0A",X"1F",X"3D",X"06",X"0C",X"03",X"0C",X"0E",X"1F",X"85",X"06",X"0C",X"03",X"0C",X"FF",X"0A",
		X"32",X"A4",X"08",X"11",X"04",X"11",X"0E",X"33",X"2C",X"08",X"11",X"04",X"11",X"FF",X"0A",X"1D",
		X"C3",X"09",X"13",X"04",X"13",X"0E",X"1E",X"6E",X"09",X"13",X"04",X"13",X"FF",X"09",X"17",X"04",
		X"16",X"4E",X"D9",X"33",X"B4",X"4D",X"E3",X"48",X"00",X"1A",X"33",X"B4",X"08",X"34",X"83",X"08",
		X"35",X"52",X"00",X"06",X"10",X"03",X"0F",X"4E",X"EF",X"36",X"21",X"4D",X"E3",X"48",X"00",X"22",
		X"36",X"21",X"08",X"36",X"81",X"08",X"36",X"E1",X"00",X"BD",X"53",X"FB",X"BD",X"3F",X"5E",X"BD",
		X"4F",X"F7",X"BD",X"3E",X"8F",X"CE",X"51",X"39",X"10",X"8E",X"B2",X"5E",X"8E",X"00",X"08",X"BD",
		X"7F",X"33",X"CC",X"00",X"00",X"97",X"39",X"97",X"D0",X"DD",X"DD",X"97",X"D3",X"97",X"D4",X"97",
		X"D1",X"97",X"D2",X"97",X"DB",X"97",X"E9",X"86",X"FF",X"97",X"52",X"86",X"0A",X"97",X"3F",X"86",
		X"80",X"D6",X"E4",X"27",X"05",X"BD",X"3E",X"23",X"86",X"01",X"97",X"43",X"B6",X"A9",X"14",X"80",
		X"05",X"97",X"F2",X"0F",X"F3",X"96",X"E3",X"81",X"0A",X"27",X"08",X"81",X"0F",X"27",X"04",X"81",
		X"10",X"26",X"02",X"03",X"F3",X"86",X"0F",X"97",X"67",X"CC",X"02",X"FE",X"97",X"ED",X"97",X"EC",
		X"D7",X"EF",X"D7",X"EE",X"0D",X"E1",X"27",X"04",X"03",X"EC",X"03",X"EF",X"96",X"E3",X"48",X"CE",
		X"54",X"5D",X"8E",X"B0",X"6C",X"AD",X"D6",X"BD",X"50",X"6E",X"BD",X"50",X"A4",X"BD",X"39",X"5D",
		X"8E",X"54",X"85",X"BD",X"50",X"4E",X"BF",X"BB",X"9F",X"FD",X"BB",X"A1",X"8E",X"54",X"85",X"BD",
		X"50",X"4E",X"BF",X"A8",X"DA",X"FD",X"A8",X"DC",X"8E",X"54",X"97",X"BD",X"50",X"4E",X"BF",X"A8",
		X"D5",X"FD",X"A8",X"D7",X"8E",X"54",X"A9",X"BD",X"50",X"4E",X"BF",X"AF",X"7A",X"FD",X"AF",X"7C",
		X"8E",X"54",X"85",X"BD",X"50",X"4E",X"BF",X"A8",X"F4",X"FD",X"A8",X"F6",X"CC",X"05",X"00",X"FD",
		X"AF",X"F7",X"CC",X"00",X"00",X"B3",X"AF",X"F7",X"FD",X"AF",X"F9",X"BD",X"50",X"2C",X"B7",X"BB",
		X"B7",X"B7",X"A8",X"F2",X"B7",X"AF",X"7E",X"B7",X"A8",X"D9",X"B7",X"A8",X"F8",X"7F",X"AF",X"FB",
		X"8E",X"54",X"BB",X"8D",X"2B",X"B7",X"BB",X"B8",X"B7",X"A8",X"F3",X"B7",X"AF",X"7F",X"B7",X"A8",
		X"F9",X"CC",X"A4",X"00",X"DD",X"D9",X"39",X"DC",X"10",X"27",X"14",X"CE",X"B1",X"FE",X"37",X"36",
		X"10",X"83",X"FF",X"FF",X"27",X"09",X"34",X"40",X"BD",X"63",X"61",X"35",X"40",X"20",X"EF",X"39",
		X"C6",X"08",X"96",X"F3",X"27",X"02",X"C6",X"06",X"96",X"E1",X"3D",X"34",X"04",X"96",X"E3",X"A6",
		X"86",X"AB",X"E0",X"9B",X"F2",X"81",X"36",X"23",X"02",X"86",X"36",X"39",X"86",X"04",X"F6",X"A9",
		X"14",X"C1",X"04",X"25",X"08",X"C1",X"06",X"23",X"0E",X"86",X"03",X"20",X"0A",X"C1",X"02",X"25",
		X"04",X"86",X"05",X"20",X"02",X"86",X"06",X"D6",X"F3",X"27",X"02",X"8B",X"01",X"39",X"96",X"E1",
		X"C6",X"40",X"3D",X"34",X"06",X"96",X"E2",X"48",X"EC",X"86",X"E3",X"E1",X"10",X"83",X"03",X"C0",
		X"23",X"03",X"CC",X"03",X"C0",X"34",X"06",X"CC",X"00",X"00",X"A3",X"E4",X"35",X"90",X"8E",X"B0",
		X"74",X"EC",X"84",X"2A",X"04",X"84",X"7F",X"A7",X"84",X"EC",X"08",X"2A",X"0C",X"10",X"83",X"FF",
		X"FF",X"27",X"20",X"84",X"7F",X"A7",X"08",X"20",X"16",X"A3",X"84",X"10",X"83",X"00",X"80",X"25",
		X"02",X"C6",X"7F",X"BD",X"3E",X"78",X"96",X"D5",X"3D",X"EE",X"84",X"33",X"C6",X"EF",X"84",X"30",
		X"08",X"20",X"D6",X"39",X"8E",X"B0",X"6C",X"EC",X"84",X"10",X"83",X"FF",X"FF",X"27",X"3F",X"A6",
		X"03",X"81",X"02",X"27",X"04",X"30",X"08",X"20",X"EE",X"BD",X"3E",X"78",X"96",X"D5",X"84",X"03",
		X"CE",X"51",X"09",X"A6",X"C6",X"A7",X"04",X"BD",X"3E",X"78",X"86",X"1E",X"D6",X"D6",X"3D",X"8B",
		X"3A",X"A7",X"06",X"96",X"E1",X"CE",X"50",X"EF",X"E6",X"C6",X"DB",X"F2",X"34",X"04",X"CE",X"50",
		X"FC",X"A6",X"C6",X"D6",X"D5",X"3D",X"AB",X"E0",X"84",X"1F",X"A7",X"07",X"20",X"C7",X"39",X"0A",
		X"0C",X"0C",X"10",X"10",X"14",X"14",X"14",X"14",X"18",X"18",X"18",X"18",X"04",X"0C",X"10",X"0C",
		X"0C",X"08",X"08",X"0A",X"0A",X"06",X"06",X"06",X"06",X"20",X"30",X"60",X"70",X"1C",X"1E",X"16",
		X"14",X"10",X"12",X"1C",X"14",X"1E",X"16",X"16",X"37",X"28",X"37",X"48",X"38",X"6D",X"37",X"85",
		X"37",X"13",X"B1",X"7E",X"B1",X"34",X"3A",X"5F",X"3A",X"01",X"CC",X"8F",X"CC",X"25",X"90",X"6D",
		X"90",X"01",X"39",X"8F",X"39",X"28",X"71",X"6C",X"71",X"02",X"04",X"08",X"0A",X"0C",X"0E",X"20",
		X"22",X"CE",X"51",X"13",X"96",X"D5",X"84",X"01",X"A6",X"C6",X"CE",X"51",X"15",X"EE",X"C6",X"EF",
		X"06",X"39",X"BD",X"3E",X"78",X"30",X"08",X"EC",X"84",X"10",X"83",X"FF",X"FF",X"39",X"CE",X"51",
		X"15",X"EE",X"C6",X"EF",X"04",X"A7",X"02",X"39",X"C6",X"03",X"8D",X"17",X"BD",X"51",X"5E",X"6F",
		X"02",X"C6",X"1E",X"A6",X"04",X"81",X"49",X"23",X"02",X"C6",X"1C",X"CE",X"51",X"15",X"EE",X"C5",
		X"EF",X"06",X"39",X"34",X"04",X"CE",X"B2",X"5E",X"D6",X"D5",X"E4",X"E4",X"A6",X"C5",X"26",X"07",
		X"BD",X"3E",X"78",X"DB",X"D6",X"20",X"F3",X"6F",X"C5",X"35",X"84",X"C6",X"07",X"8D",X"E4",X"BD",
		X"51",X"5E",X"6F",X"02",X"CE",X"51",X"15",X"E6",X"04",X"C1",X"49",X"23",X"03",X"CE",X"51",X"13",
		X"D6",X"D6",X"C4",X"01",X"E6",X"C5",X"CE",X"51",X"15",X"EE",X"C5",X"EF",X"06",X"39",X"FE",X"51",
		X"29",X"D6",X"D6",X"C4",X"01",X"27",X"03",X"FE",X"51",X"2B",X"EF",X"06",X"39",X"A6",X"02",X"81",
		X"FE",X"26",X"0C",X"96",X"D5",X"84",X"03",X"CE",X"51",X"0D",X"A6",X"C6",X"BD",X"51",X"5E",X"BD",
		X"51",X"52",X"26",X"E9",X"39",X"A6",X"03",X"81",X"20",X"26",X"03",X"BD",X"51",X"9B",X"BD",X"51",
		X"52",X"26",X"F2",X"39",X"CC",X"FF",X"FF",X"ED",X"88",X"60",X"39",X"A6",X"02",X"81",X"FE",X"26",
		X"0C",X"96",X"D5",X"84",X"01",X"CE",X"51",X"0D",X"A6",X"C6",X"BD",X"51",X"5E",X"BD",X"51",X"52",
		X"26",X"E9",X"39",X"A6",X"03",X"81",X"20",X"26",X"03",X"BD",X"51",X"41",X"BD",X"51",X"52",X"26",
		X"F2",X"39",X"CC",X"FF",X"FF",X"ED",X"88",X"58",X"A6",X"02",X"81",X"FE",X"26",X"17",X"E6",X"03",
		X"C1",X"20",X"26",X"05",X"BD",X"51",X"9B",X"20",X"0C",X"96",X"D5",X"84",X"03",X"CE",X"51",X"0D",
		X"A6",X"C6",X"BD",X"51",X"5E",X"BD",X"51",X"52",X"26",X"DE",X"39",X"A6",X"02",X"81",X"FE",X"26",
		X"0C",X"96",X"D5",X"84",X"03",X"CE",X"51",X"0D",X"A6",X"C6",X"BD",X"51",X"5E",X"BD",X"51",X"52",
		X"26",X"E9",X"39",X"A6",X"02",X"81",X"FE",X"26",X"0D",X"96",X"D5",X"C6",X"06",X"3D",X"CE",X"51",
		X"0D",X"A6",X"C6",X"BD",X"51",X"5E",X"BD",X"51",X"52",X"26",X"E8",X"8E",X"B0",X"6C",X"D6",X"E1",
		X"A6",X"03",X"81",X"04",X"26",X"07",X"5A",X"2D",X"0D",X"86",X"06",X"A7",X"03",X"34",X"04",X"BD",
		X"51",X"52",X"35",X"04",X"26",X"EA",X"39",X"81",X"01",X"23",X"04",X"86",X"20",X"A7",X"0B",X"A6",
		X"02",X"81",X"FE",X"26",X"17",X"E6",X"03",X"C1",X"20",X"26",X"05",X"BD",X"51",X"9B",X"20",X"0C",
		X"96",X"D5",X"84",X"03",X"CE",X"51",X"0D",X"A6",X"C6",X"BD",X"51",X"5E",X"BD",X"51",X"52",X"26",
		X"DE",X"39",X"96",X"E1",X"81",X"05",X"25",X"08",X"86",X"00",X"A7",X"88",X"73",X"A7",X"88",X"7B",
		X"A6",X"02",X"81",X"FE",X"26",X"17",X"E6",X"03",X"C1",X"20",X"26",X"05",X"BD",X"51",X"9B",X"20",
		X"0C",X"96",X"D5",X"84",X"01",X"CE",X"51",X"0D",X"A6",X"C6",X"BD",X"51",X"5E",X"BD",X"51",X"52",
		X"26",X"DE",X"39",X"96",X"E1",X"81",X"02",X"23",X"04",X"86",X"20",X"A7",X"0B",X"E6",X"03",X"C1",
		X"20",X"26",X"05",X"BD",X"51",X"68",X"20",X"0C",X"96",X"D5",X"84",X"01",X"CE",X"51",X"0D",X"A6",
		X"C6",X"BD",X"51",X"5E",X"BD",X"51",X"52",X"26",X"E4",X"39",X"96",X"E1",X"81",X"01",X"23",X"04",
		X"86",X"20",X"A7",X"0B",X"A6",X"02",X"81",X"FE",X"26",X"25",X"E6",X"03",X"C1",X"20",X"26",X"05",
		X"BD",X"51",X"9B",X"20",X"1A",X"96",X"D5",X"84",X"03",X"CE",X"51",X"0D",X"A6",X"C6",X"BD",X"51",
		X"5E",X"EF",X"06",X"A6",X"06",X"2B",X"04",X"86",X"10",X"20",X"02",X"86",X"80",X"A7",X"06",X"BD",
		X"51",X"52",X"26",X"D0",X"39",X"EC",X"88",X"56",X"C0",X"07",X"ED",X"06",X"96",X"E1",X"81",X"01",
		X"23",X"04",X"86",X"20",X"A7",X"0B",X"BD",X"52",X"28",X"39",X"CC",X"FF",X"FF",X"ED",X"89",X"00",
		X"88",X"A6",X"02",X"81",X"FE",X"26",X"17",X"E6",X"03",X"C1",X"20",X"26",X"05",X"BD",X"51",X"9B",
		X"20",X"0C",X"96",X"D5",X"84",X"03",X"CE",X"51",X"0D",X"A6",X"C6",X"BD",X"51",X"5E",X"BD",X"51",
		X"52",X"26",X"DE",X"39",X"96",X"D5",X"84",X"0F",X"B7",X"B2",X"5D",X"7F",X"B2",X"5C",X"CE",X"B2",
		X"3C",X"86",X"10",X"34",X"02",X"86",X"26",X"8B",X"04",X"BD",X"3E",X"78",X"D6",X"D5",X"C4",X"7F",
		X"CB",X"50",X"ED",X"C1",X"6A",X"E4",X"26",X"EF",X"35",X"02",X"A6",X"03",X"81",X"30",X"26",X"10",
		X"CE",X"B2",X"3C",X"B6",X"B2",X"5C",X"7C",X"B2",X"5C",X"48",X"EC",X"C6",X"ED",X"06",X"20",X"11",
		X"81",X"20",X"26",X"09",X"8D",X"11",X"ED",X"04",X"BD",X"51",X"BE",X"20",X"04",X"8D",X"08",X"ED",
		X"06",X"BD",X"51",X"52",X"26",X"D4",X"39",X"B6",X"B2",X"5D",X"8B",X"07",X"84",X"0F",X"B7",X"B2",
		X"5D",X"CE",X"B2",X"3C",X"48",X"EC",X"C6",X"C0",X"06",X"39",X"39",X"0F",X"E4",X"0F",X"EA",X"0F",
		X"EB",X"0F",X"E1",X"DC",X"10",X"8D",X"4A",X"D7",X"E2",X"4F",X"0D",X"E1",X"27",X"02",X"86",X"08",
		X"9B",X"E2",X"97",X"E3",X"96",X"11",X"81",X"64",X"26",X"04",X"86",X"11",X"97",X"E3",X"D6",X"E2",
		X"C1",X"08",X"26",X"02",X"03",X"E4",X"96",X"E3",X"81",X"09",X"26",X"0F",X"96",X"E1",X"84",X"01",
		X"27",X"1A",X"CC",X"FF",X"12",X"97",X"EA",X"D7",X"E3",X"20",X"11",X"81",X"0A",X"26",X"0D",X"96",
		X"E1",X"84",X"01",X"26",X"07",X"CC",X"FF",X"13",X"97",X"EB",X"D7",X"E3",X"96",X"E1",X"D6",X"E2",
		X"39",X"83",X"00",X"08",X"2F",X"04",X"0C",X"E1",X"20",X"F7",X"CB",X"08",X"39",X"51",X"CD",X"51",
		X"CD",X"51",X"E5",X"51",X"F4",X"51",X"FB",X"52",X"13",X"52",X"22",X"52",X"4B",X"52",X"63",X"52",
		X"97",X"52",X"D0",X"51",X"FA",X"52",X"F3",X"53",X"1A",X"53",X"55",X"52",X"C2",X"52",X"63",X"53",
		X"6A",X"53",X"94",X"53",X"FA",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",
		X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",X"03",
		X"80",X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",X"01",X"80",X"02",X"00",X"02",X"00",X"02",
		X"00",X"02",X"40",X"02",X"40",X"02",X"80",X"02",X"80",X"02",X"C0",X"08",X"08",X"08",X"0E",X"0E",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0C",X"0E",X"0E",X"0E",X"0E",X"0C",X"0C",X"0E",X"0E",X"0E",X"34",
		X"01",X"1A",X"50",X"C6",X"02",X"BD",X"E5",X"61",X"BD",X"E0",X"E5",X"4F",X"5F",X"FD",X"AF",X"75",
		X"CE",X"58",X"B3",X"BD",X"E4",X"20",X"BD",X"57",X"22",X"BD",X"57",X"14",X"8E",X"55",X"D0",X"BD",
		X"F4",X"44",X"8E",X"55",X"D7",X"BD",X"F4",X"44",X"8E",X"55",X"DE",X"BD",X"F4",X"44",X"8E",X"56",
		X"02",X"BD",X"F5",X"4F",X"8E",X"56",X"2F",X"BD",X"F5",X"4F",X"8E",X"56",X"54",X"BD",X"F5",X"4F",
		X"8E",X"55",X"E5",X"BD",X"F5",X"CC",X"1C",X"AF",X"BD",X"E5",X"1F",X"BD",X"57",X"6B",X"FC",X"AF",
		X"75",X"10",X"83",X"03",X"83",X"25",X"F1",X"CC",X"0C",X"A4",X"FD",X"AF",X"77",X"8D",X"39",X"DC",
		X"D5",X"84",X"07",X"8B",X"03",X"BB",X"AF",X"77",X"B7",X"AF",X"77",X"81",X"7F",X"22",X"1F",X"C4",
		X"0F",X"C0",X"0A",X"FB",X"AF",X"78",X"C1",X"1A",X"22",X"02",X"C6",X"1A",X"F7",X"AF",X"78",X"86",
		X"06",X"B7",X"AF",X"79",X"BD",X"E5",X"1F",X"7A",X"AF",X"79",X"26",X"F8",X"20",X"CF",X"86",X"78",
		X"BD",X"E5",X"1F",X"4A",X"26",X"FA",X"35",X"81",X"34",X"01",X"1A",X"50",X"86",X"01",X"BD",X"70",
		X"08",X"BD",X"00",X"A2",X"BD",X"F8",X"B5",X"CC",X"00",X"00",X"ED",X"42",X"CC",X"01",X"01",X"ED",
		X"46",X"CC",X"0A",X"00",X"ED",X"40",X"FC",X"AF",X"77",X"ED",X"44",X"86",X"05",X"A7",X"C8",X"1F",
		X"CC",X"55",X"97",X"ED",X"4A",X"35",X"81",X"6F",X"C8",X"30",X"CC",X"08",X"0E",X"ED",X"46",X"CC",
		X"55",X"A6",X"ED",X"4A",X"20",X"05",X"6A",X"C8",X"1C",X"26",X"1E",X"86",X"04",X"A7",X"C8",X"1C",
		X"6C",X"C8",X"30",X"A6",X"C8",X"30",X"81",X"04",X"25",X"05",X"BD",X"F9",X"16",X"20",X"0A",X"8E",
		X"55",X"C8",X"48",X"EC",X"86",X"ED",X"42",X"6C",X"4F",X"39",X"00",X"00",X"00",X"70",X"00",X"E0",
		X"00",X"00",X"00",X"66",X"25",X"2C",X"15",X"03",X"9C",X"00",X"34",X"44",X"5E",X"28",X"12",X"4C",
		X"00",X"3E",X"72",X"55",X"28",X"55",X"EB",X"00",X"50",X"A5",X"DD",X"54",X"48",X"45",X"20",X"44",
		X"41",X"59",X"20",X"54",X"48",X"45",X"59",X"20",X"54",X"4F",X"4F",X"4B",X"20",X"4F",X"56",X"45",
		X"52",X"FF",X"56",X"08",X"00",X"46",X"C4",X"44",X"44",X"45",X"53",X"49",X"47",X"4E",X"45",X"44",
		X"20",X"42",X"59",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",
		X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"2C",X"20",X"49",X"4E",X"43",X"2E",X"FF",X"56",
		X"35",X"00",X"56",X"CB",X"44",X"53",X"4F",X"46",X"54",X"57",X"41",X"52",X"45",X"20",X"42",X"59",
		X"20",X"47",X"41",X"4D",X"45",X"53",X"20",X"41",X"4C",X"49",X"56",X"45",X"21",X"2C",X"20",X"49",
		X"4E",X"43",X"2E",X"FF",X"56",X"5A",X"00",X"40",X"D4",X"44",X"43",X"4F",X"50",X"59",X"52",X"49",
		X"47",X"48",X"54",X"20",X"31",X"39",X"38",X"34",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",
		X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"2C",X"20",X"49",
		X"4E",X"43",X"2E",X"FF",X"F0",X"00",X"0A",X"0E",X"01",X"DC",X"D0",X"00",X"0C",X"10",X"01",X"D8",
		X"F0",X"00",X"0E",X"12",X"01",X"D4",X"D0",X"00",X"10",X"14",X"01",X"D0",X"F0",X"00",X"12",X"16",
		X"01",X"CC",X"D0",X"00",X"14",X"18",X"01",X"C8",X"0F",X"01",X"19",X"0E",X"01",X"DC",X"0D",X"01",
		X"17",X"10",X"01",X"D8",X"0F",X"01",X"15",X"12",X"01",X"D4",X"0D",X"01",X"13",X"14",X"01",X"D0",
		X"0F",X"01",X"11",X"16",X"01",X"CC",X"0D",X"01",X"0F",X"18",X"01",X"C8",X"FF",X"00",X"0A",X"0E",
		X"88",X"01",X"DD",X"00",X"0C",X"10",X"86",X"01",X"FF",X"00",X"0E",X"12",X"84",X"01",X"DD",X"00",
		X"10",X"14",X"82",X"01",X"FF",X"00",X"12",X"16",X"80",X"01",X"DD",X"00",X"14",X"18",X"7E",X"01",
		X"FF",X"00",X"0A",X"EA",X"88",X"01",X"DD",X"00",X"0C",X"E8",X"86",X"01",X"FF",X"00",X"0E",X"E6",
		X"84",X"01",X"DD",X"00",X"10",X"E4",X"82",X"01",X"FF",X"00",X"12",X"E2",X"80",X"01",X"DD",X"00",
		X"14",X"E0",X"7E",X"01",X"C6",X"18",X"8E",X"56",X"84",X"BD",X"F4",X"87",X"30",X"06",X"5A",X"26",
		X"F8",X"39",X"8E",X"AF",X"6E",X"CC",X"1F",X"42",X"ED",X"04",X"CC",X"1A",X"03",X"A7",X"03",X"F7",
		X"AF",X"74",X"CE",X"57",X"5F",X"10",X"8E",X"00",X"16",X"10",X"AF",X"01",X"86",X"04",X"E6",X"C0",
		X"E7",X"00",X"BD",X"F4",X"87",X"10",X"AE",X"01",X"31",X"A8",X"3E",X"10",X"AF",X"01",X"4A",X"26",
		X"ED",X"7A",X"AF",X"74",X"27",X"08",X"E6",X"03",X"CB",X"42",X"E7",X"03",X"20",X"D7",X"39",X"11",
		X"22",X"33",X"55",X"33",X"88",X"11",X"BB",X"22",X"BB",X"55",X"88",X"FC",X"AF",X"75",X"C3",X"00",
		X"01",X"FD",X"AF",X"75",X"CE",X"58",X"B3",X"BD",X"E3",X"EE",X"39",X"00",X"00",X"00",X"3C",X"57",
		X"81",X"4F",X"F1",X"00",X"F0",X"57",X"87",X"00",X"00",X"00",X"3C",X"57",X"8D",X"4F",X"F1",X"00",
		X"3C",X"57",X"87",X"00",X"00",X"00",X"3C",X"57",X"99",X"DF",X"F1",X"00",X"F0",X"57",X"9F",X"00",
		X"00",X"00",X"3C",X"57",X"A5",X"DF",X"F1",X"00",X"3C",X"57",X"9F",X"00",X"00",X"00",X"78",X"57",
		X"B1",X"4F",X"F1",X"00",X"B4",X"57",X"B7",X"00",X"00",X"00",X"3C",X"57",X"BD",X"4F",X"F1",X"00",
		X"3C",X"57",X"B7",X"00",X"00",X"00",X"78",X"57",X"C9",X"DF",X"F1",X"00",X"B4",X"57",X"CF",X"00",
		X"00",X"00",X"3C",X"57",X"D5",X"DF",X"F1",X"00",X"3C",X"57",X"CF",X"00",X"00",X"00",X"B4",X"57",
		X"E1",X"4F",X"F1",X"00",X"78",X"57",X"E7",X"00",X"00",X"00",X"3C",X"57",X"ED",X"4F",X"F1",X"00",
		X"3C",X"57",X"E7",X"00",X"00",X"00",X"B4",X"57",X"F9",X"DF",X"F1",X"00",X"78",X"57",X"FF",X"00",
		X"00",X"00",X"3C",X"58",X"05",X"DF",X"F1",X"00",X"3C",X"57",X"FF",X"00",X"00",X"02",X"D0",X"58",
		X"11",X"F0",X"F0",X"00",X"02",X"58",X"1D",X"00",X"00",X"02",X"D1",X"58",X"1D",X"FF",X"FF",X"00",
		X"02",X"58",X"29",X"00",X"00",X"02",X"D0",X"58",X"29",X"00",X"FF",X"00",X"02",X"58",X"35",X"00",
		X"00",X"02",X"D1",X"58",X"35",X"FF",X"F0",X"00",X"02",X"58",X"41",X"00",X"00",X"02",X"D0",X"58",
		X"41",X"F0",X"FF",X"00",X"02",X"58",X"4D",X"00",X"00",X"02",X"D1",X"58",X"4D",X"0F",X"FF",X"00",
		X"02",X"58",X"11",X"0F",X"48",X"00",X"04",X"58",X"59",X"0F",X"58",X"00",X"04",X"58",X"5F",X"0F",
		X"68",X"00",X"04",X"58",X"65",X"0F",X"78",X"00",X"04",X"58",X"6B",X"0F",X"88",X"00",X"04",X"58",
		X"71",X"0F",X"98",X"00",X"04",X"58",X"77",X"0F",X"A8",X"00",X"04",X"58",X"7D",X"0F",X"B8",X"00",
		X"04",X"58",X"83",X"0F",X"C8",X"00",X"04",X"58",X"89",X"0F",X"D8",X"00",X"04",X"58",X"8F",X"0F",
		X"E8",X"00",X"04",X"58",X"95",X"0F",X"F8",X"00",X"04",X"58",X"8F",X"0F",X"F8",X"00",X"06",X"58",
		X"A1",X"E6",X"FF",X"00",X"06",X"58",X"9B",X"E6",X"FF",X"00",X"06",X"58",X"AD",X"0F",X"F8",X"00",
		X"06",X"58",X"A7",X"0A",X"57",X"7B",X"0C",X"57",X"93",X"07",X"57",X"AB",X"09",X"57",X"C3",X"06",
		X"57",X"DB",X"0E",X"57",X"F3",X"01",X"58",X"0B",X"02",X"58",X"17",X"03",X"58",X"23",X"05",X"58",
		X"2F",X"08",X"58",X"3B",X"0B",X"58",X"47",X"04",X"58",X"53",X"0F",X"58",X"A7",X"0D",X"58",X"9B",
		X"FF",X"E6",X"C8",X"15",X"86",X"07",X"3D",X"8E",X"5B",X"1B",X"3A",X"EC",X"00",X"ED",X"C8",X"36",
		X"EC",X"02",X"ED",X"C8",X"3B",X"EC",X"04",X"ED",X"C8",X"48",X"E6",X"06",X"A6",X"C8",X"14",X"A0",
		X"C8",X"30",X"25",X"10",X"8E",X"5A",X"E4",X"3D",X"44",X"56",X"44",X"56",X"44",X"56",X"44",X"56",
		X"44",X"56",X"20",X"14",X"8E",X"5A",X"AD",X"40",X"3D",X"44",X"56",X"44",X"56",X"44",X"56",X"44",
		X"56",X"44",X"56",X"43",X"53",X"C3",X"00",X"01",X"ED",X"C8",X"34",X"AF",X"C8",X"39",X"6F",X"C8",
		X"42",X"6F",X"4E",X"6F",X"C8",X"4A",X"CC",X"FA",X"00",X"ED",X"C8",X"32",X"8E",X"59",X"F4",X"AF",
		X"C8",X"46",X"8E",X"59",X"58",X"AF",X"4A",X"C6",X"05",X"E7",X"C8",X"1F",X"A6",X"C8",X"30",X"E6",
		X"C8",X"32",X"83",X"05",X"0D",X"ED",X"44",X"39",X"96",X"40",X"26",X"07",X"A6",X"4E",X"27",X"04",
		X"BD",X"30",X"7C",X"39",X"96",X"39",X"26",X"0D",X"EC",X"C8",X"48",X"83",X"00",X"01",X"ED",X"C8",
		X"48",X"10",X"27",X"00",X"D0",X"6A",X"C8",X"42",X"2E",X"36",X"AE",X"C8",X"39",X"A6",X"80",X"26",
		X"23",X"AD",X"D8",X"46",X"27",X"0F",X"EC",X"02",X"ED",X"46",X"EC",X"04",X"ED",X"C8",X"3D",X"A6",
		X"06",X"30",X"07",X"20",X"0F",X"EC",X"84",X"ED",X"C8",X"39",X"A6",X"C8",X"4A",X"27",X"03",X"BD",
		X"70",X"08",X"20",X"0C",X"A7",X"C8",X"42",X"EC",X"81",X"ED",X"42",X"AF",X"C8",X"39",X"6C",X"4F",
		X"96",X"39",X"26",X"3F",X"EC",X"C8",X"37",X"A3",X"C8",X"3B",X"ED",X"C8",X"37",X"A6",X"C8",X"36",
		X"82",X"00",X"A7",X"C8",X"36",X"EC",X"C8",X"32",X"A3",X"C8",X"36",X"ED",X"C8",X"32",X"EC",X"C8",
		X"30",X"E3",X"C8",X"34",X"ED",X"C8",X"30",X"E6",X"C8",X"32",X"A3",X"C8",X"3D",X"10",X"A3",X"44",
		X"27",X"11",X"6C",X"4F",X"ED",X"44",X"A6",X"40",X"84",X"DF",X"E6",X"C8",X"31",X"2A",X"02",X"8A",
		X"20",X"A7",X"40",X"39",X"CC",X"59",X"FB",X"ED",X"C8",X"46",X"39",X"A6",X"C8",X"32",X"81",X"64",
		X"22",X"0C",X"CC",X"5A",X"10",X"ED",X"C8",X"46",X"86",X"13",X"A7",X"C8",X"4A",X"39",X"4F",X"39",
		X"A6",X"C8",X"32",X"81",X"1C",X"22",X"18",X"CC",X"5A",X"31",X"ED",X"C8",X"46",X"34",X"10",X"96",
		X"E4",X"26",X"05",X"86",X"03",X"BD",X"D0",X"5E",X"86",X"14",X"A7",X"C8",X"4A",X"35",X"90",X"4F",
		X"39",X"A6",X"C8",X"36",X"2B",X"02",X"4F",X"39",X"86",X"3C",X"97",X"5C",X"CC",X"5A",X"43",X"ED",
		X"C8",X"46",X"39",X"4F",X"39",X"96",X"E4",X"26",X"4A",X"8E",X"5A",X"9F",X"A6",X"C8",X"34",X"2B",
		X"03",X"8E",X"5A",X"A6",X"96",X"67",X"A7",X"4D",X"A6",X"C8",X"30",X"E6",X"C8",X"32",X"A3",X"05",
		X"ED",X"44",X"EC",X"03",X"ED",X"46",X"EC",X"01",X"ED",X"42",X"8E",X"5A",X"72",X"AF",X"4A",X"6C",
		X"4F",X"39",X"96",X"39",X"26",X"21",X"96",X"E4",X"26",X"19",X"6A",X"4D",X"2A",X"19",X"BE",X"B0",
		X"55",X"27",X"10",X"6C",X"0E",X"8E",X"31",X"FD",X"AF",X"4A",X"8E",X"42",X"86",X"AF",X"C8",X"39",
		X"6C",X"4E",X"39",X"AD",X"D8",X"22",X"39",X"A6",X"4E",X"27",X"03",X"BD",X"30",X"7C",X"39",X"14",
		X"25",X"14",X"06",X"0A",X"03",X"05",X"14",X"1B",X"5D",X"06",X"0A",X"03",X"05",X"00",X"00",X"00",
		X"0B",X"1A",X"05",X"0D",X"02",X"20",X"2D",X"00",X"5A",X"B4",X"0D",X"13",X"06",X"09",X"04",X"21",
		X"4B",X"04",X"22",X"42",X"04",X"23",X"39",X"00",X"5A",X"BE",X"06",X"0E",X"03",X"07",X"04",X"24",
		X"30",X"04",X"24",X"84",X"00",X"5A",X"CE",X"06",X"0A",X"03",X"05",X"04",X"24",X"D8",X"04",X"25",
		X"14",X"00",X"5A",X"DB",X"00",X"00",X"00",X"0B",X"1A",X"05",X"0D",X"02",X"16",X"76",X"00",X"5A",
		X"EB",X"0D",X"13",X"06",X"09",X"04",X"17",X"94",X"04",X"18",X"8B",X"04",X"19",X"82",X"00",X"5A",
		X"F5",X"06",X"0E",X"03",X"07",X"04",X"1A",X"79",X"04",X"1A",X"CD",X"00",X"5B",X"05",X"06",X"0A",
		X"03",X"05",X"04",X"1B",X"21",X"04",X"1B",X"5D",X"00",X"5B",X"12",X"02",X"AB",X"03",X"F1",X"00",
		X"CD",X"27",X"02",X"BC",X"04",X"24",X"00",X"C8",X"28",X"02",X"CF",X"04",X"5C",X"00",X"C3",X"2A",
		X"02",X"E1",X"04",X"97",X"00",X"BE",X"2B",X"02",X"F5",X"04",X"D8",X"00",X"B9",X"2C",X"03",X"0A",
		X"05",X"1D",X"00",X"B4",X"2D",X"03",X"21",X"05",X"69",X"00",X"AF",X"2E",X"03",X"39",X"05",X"BC",
		X"00",X"AA",X"30",X"03",X"52",X"06",X"16",X"00",X"A5",X"31",X"03",X"6C",X"06",X"79",X"00",X"A0",
		X"33",X"03",X"89",X"06",X"E6",X"00",X"9B",X"34",X"03",X"A7",X"07",X"5E",X"00",X"96",X"36",X"03",
		X"C7",X"07",X"E2",X"00",X"91",X"38",X"03",X"EA",X"08",X"75",X"00",X"8C",X"3A",X"04",X"10",X"09",
		X"18",X"00",X"87",X"3C",X"04",X"38",X"09",X"CF",X"00",X"82",X"3F",X"04",X"63",X"0A",X"9C",X"00",
		X"7D",X"41",X"04",X"92",X"0B",X"83",X"00",X"78",X"44",X"04",X"C6",X"0C",X"89",X"00",X"73",X"47",
		X"04",X"FD",X"0D",X"B3",X"00",X"6E",X"4A",X"05",X"3A",X"0F",X"09",X"00",X"69",X"4E",X"05",X"7D",
		X"10",X"93",X"00",X"64",X"51",X"05",X"C8",X"12",X"5E",X"00",X"5F",X"56",X"06",X"1B",X"14",X"77",
		X"00",X"5A",X"5B",X"06",X"78",X"16",X"F2",X"00",X"55",X"60",X"06",X"DF",X"19",X"E7",X"00",X"50",
		X"66",X"07",X"56",X"1D",X"78",X"00",X"4B",X"6D",X"07",X"DC",X"21",X"D5",X"00",X"46",X"75",X"08",
		X"79",X"27",X"3C",X"00",X"41",X"7E",X"09",X"30",X"2E",X"0C",X"00",X"3C",X"88",X"0A",X"08",X"36",
		X"CD",X"00",X"37",X"94",X"0B",X"0B",X"42",X"4F",X"00",X"32",X"A3",X"86",X"01",X"A7",X"C8",X"1F",
		X"F6",X"B0",X"40",X"96",X"D5",X"3D",X"BE",X"B0",X"41",X"4A",X"2B",X"05",X"AE",X"88",X"1A",X"20",
		X"F8",X"AF",X"C8",X"54",X"CC",X"30",X"44",X"ED",X"42",X"CC",X"07",X"16",X"ED",X"46",X"44",X"40",
		X"AB",X"C8",X"30",X"54",X"50",X"EB",X"C8",X"32",X"ED",X"44",X"CC",X"00",X"00",X"ED",X"C8",X"47",
		X"A7",X"4E",X"A7",X"C8",X"1D",X"ED",X"C8",X"34",X"ED",X"C8",X"36",X"A7",X"C8",X"38",X"A7",X"C8",
		X"44",X"A7",X"C8",X"45",X"A7",X"C8",X"4A",X"B6",X"AF",X"7E",X"A7",X"C8",X"3C",X"A7",X"C8",X"3B",
		X"8E",X"5C",X"67",X"AF",X"C8",X"3E",X"8E",X"5C",X"5C",X"AF",X"4A",X"39",X"A6",X"4E",X"27",X"04",
		X"BD",X"30",X"7C",X"39",X"6E",X"D8",X"3E",X"8E",X"5C",X"B6",X"AF",X"C8",X"3E",X"EC",X"C8",X"14",
		X"ED",X"C8",X"5E",X"A1",X"C8",X"30",X"25",X"19",X"22",X"1C",X"8E",X"00",X"00",X"E1",X"C8",X"32",
		X"26",X"17",X"A6",X"C8",X"1D",X"26",X"2C",X"86",X"FF",X"A7",X"C8",X"1D",X"BD",X"39",X"13",X"20",
		X"0F",X"BE",X"AF",X"7C",X"20",X"03",X"BE",X"AF",X"7A",X"E1",X"C8",X"32",X"25",X"07",X"22",X"0A",
		X"CC",X"00",X"00",X"20",X"08",X"FC",X"AF",X"7C",X"20",X"03",X"FC",X"AF",X"7A",X"ED",X"C8",X"36",
		X"AF",X"C8",X"34",X"7E",X"5E",X"AF",X"8E",X"5D",X"D4",X"AF",X"C8",X"3E",X"A6",X"C8",X"30",X"E6",
		X"C8",X"32",X"BD",X"67",X"5E",X"A7",X"C8",X"38",X"27",X"08",X"A7",X"C8",X"16",X"8E",X"5C",X"D5",
		X"AF",X"4A",X"7E",X"5E",X"AF",X"A6",X"C8",X"16",X"8E",X"5E",X"BA",X"AE",X"86",X"A6",X"C8",X"30",
		X"E6",X"C8",X"32",X"6E",X"84",X"10",X"A3",X"C8",X"5E",X"27",X"08",X"20",X"12",X"10",X"A3",X"C8",
		X"5E",X"26",X"14",X"BD",X"F9",X"16",X"39",X"C1",X"EC",X"25",X"5D",X"C6",X"EC",X"20",X"3F",X"C1",
		X"B1",X"22",X"55",X"C6",X"B1",X"20",X"27",X"C1",X"39",X"25",X"04",X"C6",X"39",X"20",X"2F",X"C1",
		X"37",X"22",X"45",X"C6",X"37",X"20",X"17",X"C1",X"38",X"22",X"3D",X"C6",X"38",X"20",X"0F",X"C1",
		X"97",X"22",X"35",X"C6",X"98",X"8E",X"00",X"00",X"AF",X"C8",X"34",X"BD",X"39",X"2F",X"E7",X"C8",
		X"32",X"EC",X"C8",X"36",X"2A",X"22",X"CC",X"00",X"00",X"ED",X"C8",X"36",X"20",X"1A",X"E7",X"C8",
		X"32",X"EC",X"C8",X"36",X"2F",X"12",X"20",X"EE",X"C1",X"68",X"25",X"0C",X"C6",X"68",X"20",X"EE",
		X"C1",X"48",X"25",X"04",X"C6",X"48",X"20",X"E6",X"CC",X"5C",X"5C",X"ED",X"4A",X"39",X"A7",X"C8",
		X"30",X"EC",X"C8",X"34",X"2A",X"F2",X"CC",X"00",X"00",X"ED",X"C8",X"34",X"20",X"EA",X"A7",X"C8",
		X"30",X"EC",X"C8",X"34",X"2F",X"E2",X"20",X"EE",X"81",X"24",X"22",X"DC",X"86",X"24",X"20",X"DE",
		X"81",X"6E",X"25",X"D4",X"86",X"6E",X"20",X"E6",X"81",X"1E",X"22",X"CC",X"86",X"1E",X"20",X"CE",
		X"81",X"75",X"25",X"C4",X"86",X"75",X"20",X"D6",X"81",X"26",X"22",X"BC",X"86",X"26",X"20",X"BE",
		X"81",X"6D",X"25",X"B4",X"86",X"6D",X"20",X"C6",X"81",X"28",X"22",X"AC",X"86",X"28",X"20",X"AE",
		X"81",X"6B",X"25",X"A4",X"86",X"6B",X"20",X"B6",X"C6",X"10",X"E7",X"C8",X"14",X"E6",X"C8",X"32",
		X"E7",X"C8",X"15",X"86",X"01",X"20",X"97",X"C6",X"80",X"E7",X"C8",X"14",X"E6",X"C8",X"32",X"E7",
		X"C8",X"15",X"20",X"9A",X"8E",X"5E",X"4F",X"AF",X"C8",X"3E",X"A6",X"C8",X"48",X"BB",X"AF",X"7F",
		X"A7",X"C8",X"48",X"24",X"0B",X"6C",X"C8",X"47",X"6A",X"C8",X"3C",X"2A",X"03",X"6F",X"C8",X"3C",
		X"EC",X"C8",X"36",X"2D",X"23",X"26",X"17",X"EC",X"C8",X"34",X"26",X"2A",X"6C",X"C8",X"4A",X"A6",
		X"C8",X"4A",X"81",X"08",X"25",X"46",X"BD",X"39",X"2F",X"6F",X"C8",X"4A",X"20",X"3E",X"E3",X"C8",
		X"32",X"A1",X"C8",X"5F",X"22",X"0A",X"20",X"0B",X"E3",X"C8",X"32",X"A1",X"C8",X"5F",X"24",X"03",
		X"A6",X"C8",X"5F",X"ED",X"C8",X"32",X"6F",X"C8",X"4A",X"EC",X"C8",X"34",X"2D",X"0C",X"27",X"1C",
		X"E3",X"C8",X"30",X"A1",X"C8",X"5E",X"22",X"0E",X"20",X"0F",X"E3",X"C8",X"30",X"A1",X"C8",X"5E",
		X"25",X"04",X"81",X"F0",X"25",X"03",X"A6",X"C8",X"5E",X"ED",X"C8",X"30",X"7E",X"5E",X"AF",X"8E",
		X"5E",X"A1",X"AF",X"C8",X"3E",X"EC",X"C8",X"34",X"2D",X"13",X"A6",X"C8",X"45",X"8B",X"FE",X"2A",
		X"02",X"86",X"04",X"A7",X"C8",X"45",X"8E",X"5E",X"B0",X"EC",X"86",X"20",X"11",X"A6",X"C8",X"45",
		X"8B",X"FE",X"2A",X"02",X"86",X"04",X"A7",X"C8",X"45",X"8E",X"5E",X"B6",X"EC",X"86",X"ED",X"42",
		X"86",X"07",X"44",X"40",X"AB",X"C8",X"30",X"A7",X"44",X"86",X"2A",X"E6",X"C8",X"31",X"2D",X"02",
		X"86",X"0A",X"A7",X"40",X"86",X"16",X"44",X"40",X"AB",X"C8",X"32",X"A7",X"45",X"6C",X"4F",X"20",
		X"0E",X"6A",X"C8",X"3B",X"2A",X"09",X"A6",X"C8",X"3C",X"A7",X"C8",X"3B",X"7E",X"5C",X"67",X"39",
		X"30",X"DE",X"30",X"44",X"2F",X"AA",X"32",X"AC",X"32",X"12",X"31",X"78",X"5D",X"07",X"5D",X"0F",
		X"5D",X"17",X"5D",X"0F",X"5D",X"07",X"5C",X"FF",X"5C",X"FF",X"5D",X"17",X"5D",X"17",X"5C",X"E5",
		X"5C",X"E5",X"5D",X"98",X"5D",X"A0",X"5C",X"ED",X"5C",X"ED",X"5D",X"A8",X"5D",X"B0",X"5C",X"F7",
		X"5D",X"88",X"5D",X"90",X"5D",X"07",X"5D",X"17",X"5D",X"0F",X"5D",X"78",X"5D",X"80",X"5C",X"FF",
		X"5D",X"1F",X"5D",X"48",X"5D",X"50",X"5D",X"B8",X"5D",X"C7",X"86",X"01",X"A7",X"C8",X"1F",X"86",
		X"FF",X"A7",X"C8",X"3B",X"CC",X"00",X"00",X"A7",X"4E",X"A7",X"C8",X"38",X"A7",X"C8",X"42",X"ED",
		X"C8",X"54",X"A7",X"C8",X"56",X"ED",X"C8",X"36",X"A7",X"C8",X"39",X"A7",X"C8",X"50",X"A7",X"C8",
		X"4F",X"A7",X"C8",X"3C",X"A7",X"C8",X"3D",X"ED",X"C8",X"3E",X"A7",X"C8",X"41",X"A7",X"C8",X"40",
		X"A6",X"C8",X"32",X"81",X"A0",X"22",X"08",X"81",X"58",X"22",X"07",X"86",X"04",X"20",X"05",X"4F",
		X"20",X"02",X"86",X"02",X"A7",X"C8",X"3A",X"8E",X"5F",X"B0",X"96",X"EA",X"27",X"05",X"8E",X"5F",
		X"92",X"20",X"07",X"96",X"EB",X"27",X"03",X"8E",X"5F",X"75",X"AF",X"C8",X"34",X"8E",X"5F",X"6A",
		X"96",X"E4",X"27",X"03",X"8E",X"5F",X"69",X"AF",X"4A",X"39",X"A6",X"C8",X"50",X"27",X"03",X"7E",
		X"61",X"EC",X"6E",X"D8",X"34",X"BE",X"B0",X"55",X"A6",X"88",X"32",X"A1",X"C8",X"32",X"27",X"03",
		X"AE",X"88",X"1A",X"A6",X"88",X"30",X"A1",X"C8",X"30",X"25",X"06",X"8E",X"61",X"01",X"AF",X"C8",
		X"34",X"39",X"8D",X"31",X"A6",X"C8",X"41",X"26",X"10",X"A6",X"C8",X"3D",X"27",X"11",X"AE",X"C8",
		X"3E",X"27",X"0C",X"CC",X"00",X"00",X"ED",X"88",X"3E",X"8E",X"61",X"10",X"AF",X"C8",X"34",X"39",
		X"A6",X"C8",X"42",X"27",X"0D",X"6A",X"C8",X"42",X"26",X"0A",X"8E",X"60",X"7B",X"AF",X"C8",X"34",
		X"20",X"02",X"8D",X"01",X"39",X"AE",X"C8",X"54",X"27",X"07",X"A6",X"88",X"56",X"2B",X"02",X"20",
		X"0F",X"8D",X"25",X"AF",X"C8",X"54",X"27",X"1F",X"86",X"01",X"A7",X"88",X"56",X"6F",X"C8",X"56",
		X"11",X"A3",X"88",X"54",X"26",X"11",X"A6",X"88",X"1E",X"26",X"0C",X"6F",X"88",X"1D",X"A6",X"C8",
		X"30",X"E6",X"C8",X"32",X"ED",X"88",X"14",X"39",X"86",X"FF",X"B7",X"AF",X"80",X"B7",X"AF",X"81",
		X"BE",X"B0",X"09",X"27",X"17",X"A6",X"0E",X"26",X"0E",X"A6",X"06",X"81",X"01",X"27",X"08",X"11",
		X"A3",X"88",X"54",X"26",X"02",X"8D",X"3B",X"AE",X"88",X"1A",X"26",X"E9",X"BE",X"B0",X"0D",X"27",
		X"17",X"A6",X"0E",X"26",X"0E",X"A6",X"06",X"81",X"01",X"27",X"08",X"11",X"A3",X"88",X"54",X"26",
		X"02",X"8D",X"1F",X"AE",X"88",X"1A",X"26",X"E9",X"B6",X"AF",X"80",X"81",X"FF",X"26",X"05",X"8E",
		X"00",X"00",X"20",X"0D",X"B1",X"AF",X"81",X"22",X"05",X"BE",X"AF",X"82",X"20",X"03",X"BE",X"AF",
		X"84",X"39",X"A6",X"88",X"30",X"A0",X"C8",X"30",X"2A",X"01",X"40",X"B1",X"AF",X"80",X"24",X"06",
		X"B7",X"AF",X"80",X"BF",X"AF",X"82",X"A6",X"88",X"32",X"A0",X"C8",X"32",X"2A",X"01",X"40",X"B1",
		X"AF",X"81",X"24",X"06",X"B7",X"AF",X"81",X"BF",X"AF",X"84",X"39",X"6F",X"4E",X"8E",X"60",X"83",
		X"AF",X"C8",X"34",X"AE",X"C8",X"54",X"27",X"0B",X"A6",X"0E",X"26",X"04",X"A6",X"4E",X"27",X"0E",
		X"6F",X"88",X"56",X"6F",X"C8",X"56",X"8E",X"61",X"10",X"AF",X"C8",X"34",X"20",X"40",X"BD",X"5F",
		X"F8",X"AF",X"C8",X"36",X"27",X"2E",X"EC",X"04",X"A0",X"44",X"2A",X"01",X"40",X"81",X"04",X"22",
		X"23",X"E0",X"45",X"2A",X"01",X"50",X"C1",X"04",X"22",X"1A",X"96",X"D6",X"81",X"C0",X"25",X"14",
		X"A6",X"88",X"1E",X"26",X"0F",X"10",X"AE",X"C8",X"54",X"6F",X"A8",X"56",X"86",X"FF",X"A7",X"88",
		X"56",X"AF",X"C8",X"54",X"8D",X"0B",X"E6",X"88",X"32",X"CB",X"FE",X"E7",X"C8",X"32",X"7E",X"62",
		X"D8",X"A6",X"C8",X"56",X"2A",X"1A",X"AE",X"C8",X"54",X"E6",X"88",X"30",X"A6",X"88",X"34",X"2D",
		X"06",X"2E",X"08",X"CB",X"00",X"20",X"06",X"C0",X"03",X"20",X"02",X"CB",X"00",X"E7",X"C8",X"30",
		X"39",X"96",X"D5",X"C6",X"0C",X"3D",X"8B",X"20",X"A7",X"C8",X"39",X"8E",X"61",X"1E",X"20",X"08",
		X"86",X"08",X"A7",X"C8",X"39",X"8E",X"61",X"27",X"AF",X"C8",X"34",X"7E",X"62",X"D8",X"EC",X"C8",
		X"30",X"C3",X"00",X"80",X"ED",X"C8",X"30",X"A6",X"C8",X"3A",X"A7",X"C8",X"3B",X"A6",X"C8",X"39",
		X"4A",X"2D",X"08",X"A7",X"C8",X"39",X"6C",X"C8",X"32",X"20",X"37",X"86",X"02",X"A7",X"C8",X"38",
		X"A6",X"C8",X"32",X"80",X"03",X"A7",X"C8",X"32",X"8E",X"00",X"00",X"AF",X"C8",X"54",X"6F",X"C8",
		X"56",X"D6",X"D4",X"27",X"17",X"BD",X"26",X"4F",X"C0",X"04",X"1F",X"01",X"80",X"03",X"1F",X"02",
		X"4F",X"D6",X"D4",X"34",X"40",X"BD",X"63",X"61",X"35",X"40",X"0F",X"D4",X"8E",X"61",X"75",X"AF",
		X"C8",X"34",X"7E",X"62",X"D8",X"BD",X"5F",X"C5",X"AE",X"C8",X"54",X"27",X"2D",X"A6",X"88",X"30",
		X"A0",X"C8",X"30",X"2A",X"01",X"40",X"81",X"07",X"22",X"20",X"A6",X"88",X"32",X"A0",X"C8",X"32",
		X"2A",X"01",X"40",X"81",X"07",X"22",X"13",X"A6",X"88",X"1E",X"26",X"0E",X"86",X"FF",X"A7",X"C8",
		X"56",X"A7",X"88",X"56",X"8E",X"61",X"AD",X"AF",X"C8",X"34",X"7E",X"62",X"D8",X"6F",X"C8",X"38",
		X"86",X"05",X"A7",X"C8",X"39",X"8E",X"61",X"BE",X"AF",X"C8",X"34",X"7E",X"62",X"D8",X"A6",X"C8",
		X"3A",X"A7",X"C8",X"3B",X"A6",X"C8",X"39",X"4A",X"2D",X"0B",X"A7",X"C8",X"39",X"6A",X"C8",X"32",
		X"BD",X"60",X"E1",X"20",X"14",X"AE",X"C8",X"54",X"27",X"09",X"EC",X"C8",X"14",X"ED",X"88",X"14",
		X"6F",X"88",X"1D",X"8E",X"60",X"7B",X"AF",X"C8",X"34",X"7E",X"62",X"D8",X"6F",X"C8",X"50",X"86",
		X"08",X"A7",X"C8",X"1C",X"CC",X"01",X"01",X"ED",X"46",X"8E",X"62",X"01",X"AF",X"C8",X"34",X"20",
		X"0D",X"6A",X"C8",X"1C",X"26",X"06",X"8E",X"62",X"22",X"AF",X"C8",X"34",X"8D",X"01",X"39",X"BD",
		X"26",X"4F",X"80",X"01",X"CB",X"03",X"A7",X"C8",X"30",X"E7",X"C8",X"32",X"C0",X"0A",X"ED",X"C8",
		X"14",X"39",X"8E",X"70",X"C1",X"BD",X"6F",X"D3",X"86",X"1E",X"A7",X"C8",X"1C",X"6F",X"4E",X"96",
		X"98",X"2A",X"08",X"8E",X"01",X"91",X"CC",X"07",X"0E",X"20",X"06",X"8E",X"00",X"ED",X"CC",X"07",
		X"0E",X"AF",X"42",X"ED",X"46",X"8E",X"62",X"4B",X"AF",X"C8",X"34",X"A6",X"C8",X"1C",X"27",X"08",
		X"6A",X"C8",X"1C",X"26",X"03",X"BD",X"25",X"F9",X"8D",X"B5",X"8D",X"19",X"6C",X"4F",X"8D",X"33",
		X"A6",X"4E",X"27",X"0E",X"8E",X"61",X"10",X"AF",X"C8",X"34",X"BD",X"26",X"2C",X"C0",X"07",X"ED",
		X"C8",X"14",X"7E",X"63",X"14",X"A6",X"46",X"44",X"40",X"AB",X"C8",X"30",X"A7",X"44",X"86",X"2A",
		X"E6",X"C8",X"31",X"2D",X"02",X"86",X"0A",X"A7",X"40",X"A6",X"47",X"44",X"40",X"AB",X"C8",X"32",
		X"A7",X"45",X"39",X"34",X"02",X"E6",X"C8",X"30",X"C1",X"F0",X"25",X"04",X"C6",X"03",X"20",X"19",
		X"C1",X"20",X"22",X"04",X"8D",X"21",X"20",X"1D",X"C1",X"70",X"24",X"05",X"6F",X"C8",X"3C",X"20",
		X"14",X"8D",X"14",X"C1",X"8F",X"25",X"0E",X"C6",X"8F",X"E7",X"C8",X"30",X"8D",X"B7",X"6C",X"4F",
		X"C6",X"FE",X"E7",X"C8",X"40",X"35",X"82",X"A6",X"C8",X"3C",X"26",X"0B",X"8E",X"70",X"79",X"BD",
		X"6F",X"D3",X"86",X"FF",X"A7",X"C8",X"3C",X"39",X"A6",X"C8",X"3B",X"2D",X"45",X"A7",X"C8",X"3A",
		X"C6",X"FF",X"E7",X"C8",X"3B",X"8D",X"AC",X"A6",X"C8",X"3A",X"48",X"AB",X"C8",X"38",X"8E",X"63",
		X"49",X"AE",X"86",X"AF",X"42",X"E6",X"C8",X"56",X"2A",X"0E",X"AE",X"C8",X"54",X"AE",X"06",X"8C",
		X"01",X"01",X"26",X"04",X"AF",X"46",X"20",X"0A",X"8E",X"63",X"55",X"EC",X"86",X"ED",X"46",X"BD",
		X"62",X"75",X"6C",X"4F",X"A6",X"C8",X"40",X"81",X"FE",X"26",X"07",X"97",X"40",X"A7",X"4E",X"BD",
		X"30",X"7C",X"39",X"BE",X"B0",X"41",X"27",X"20",X"86",X"FF",X"B7",X"AF",X"80",X"B7",X"AF",X"81",
		X"BD",X"60",X"52",X"AE",X"88",X"1A",X"26",X"F8",X"B6",X"AF",X"80",X"B1",X"AF",X"81",X"22",X"05",
		X"BE",X"AF",X"82",X"20",X"03",X"BE",X"AF",X"84",X"39",X"02",X"35",X"03",X"5B",X"02",X"BA",X"03",
		X"E0",X"03",X"1A",X"04",X"40",X"07",X"13",X"07",X"13",X"06",X"10",X"06",X"10",X"05",X"0D",X"05",
		X"0D",X"34",X"01",X"1A",X"50",X"5D",X"27",X"48",X"CE",X"65",X"69",X"AD",X"D5",X"26",X"41",X"A7",
		X"C8",X"17",X"E7",X"4C",X"A6",X"4C",X"44",X"8B",X"1F",X"BD",X"70",X"08",X"1F",X"10",X"E7",X"C8",
		X"32",X"6F",X"C8",X"33",X"5F",X"ED",X"C8",X"30",X"10",X"AF",X"C8",X"14",X"6F",X"C8",X"1E",X"6F",
		X"C8",X"27",X"8E",X"67",X"B5",X"AF",X"42",X"8E",X"01",X"01",X"AF",X"46",X"8E",X"0A",X"00",X"AF",
		X"40",X"86",X"01",X"A7",X"C8",X"1F",X"A6",X"C8",X"17",X"8E",X"64",X"B0",X"AE",X"86",X"AF",X"4A",
		X"35",X"81",X"34",X"01",X"1A",X"50",X"20",X"B7",X"CC",X"14",X"30",X"20",X"12",X"CC",X"26",X"30",
		X"20",X"0D",X"CC",X"46",X"30",X"20",X"08",X"CC",X"6B",X"30",X"20",X"03",X"CC",X"83",X"30",X"8E",
		X"64",X"F0",X"20",X"73",X"CC",X"10",X"A1",X"8E",X"64",X"FE",X"20",X"6B",X"CC",X"7D",X"A1",X"8E",
		X"65",X"05",X"20",X"63",X"CC",X"31",X"31",X"8E",X"65",X"28",X"20",X"5B",X"CC",X"5C",X"31",X"8E",
		X"65",X"36",X"20",X"53",X"6A",X"C8",X"1C",X"26",X"63",X"8E",X"64",X"F7",X"20",X"4B",X"6A",X"C8",
		X"1C",X"26",X"59",X"8E",X"65",X"05",X"20",X"41",X"6A",X"C8",X"1C",X"26",X"4F",X"8E",X"65",X"0C",
		X"20",X"37",X"6A",X"C8",X"1C",X"26",X"45",X"8E",X"65",X"1A",X"20",X"2D",X"6A",X"C8",X"1C",X"26",
		X"3B",X"8E",X"65",X"21",X"20",X"23",X"8E",X"64",X"DB",X"20",X"03",X"8E",X"64",X"E9",X"A6",X"C8",
		X"30",X"80",X"05",X"20",X"0B",X"8E",X"64",X"D4",X"20",X"03",X"8E",X"64",X"E2",X"A6",X"C8",X"30",
		X"C6",X"16",X"54",X"50",X"EB",X"C8",X"32",X"ED",X"44",X"A6",X"80",X"A7",X"C8",X"1C",X"EC",X"81",
		X"ED",X"42",X"EC",X"81",X"ED",X"46",X"EC",X"84",X"ED",X"4A",X"6C",X"4F",X"39",X"E6",X"4C",X"8E",
		X"64",X"7A",X"AE",X"85",X"AF",X"4A",X"20",X"F2",X"6A",X"C8",X"1C",X"26",X"EF",X"8E",X"65",X"2F",
		X"20",X"D7",X"6A",X"C8",X"1C",X"26",X"E5",X"8E",X"65",X"3D",X"20",X"CD",X"58",X"E1",X"72",X"7B",
		X"14",X"0F",X"2B",X"BB",X"5B",X"FB",X"1B",X"52",X"69",X"C6",X"1F",X"F1",X"4D",X"30",X"00",X"00",
		X"00",X"00",X"24",X"55",X"24",X"45",X"24",X"37",X"00",X"00",X"5E",X"FA",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"47",X"C9",X"3D",X"07",X"4D",X"1F",X"4D",X"41",X"D0",X"79",X"00",X"00",
		X"64",X"5D",X"63",X"B8",X"63",X"BD",X"63",X"C2",X"63",X"C7",X"63",X"CC",X"63",X"D4",X"63",X"DC",
		X"63",X"E4",X"63",X"EC",X"64",X"5D",X"64",X"5D",X"64",X"26",X"64",X"35",X"64",X"5D",X"64",X"5D",
		X"64",X"2B",X"64",X"3A",X"08",X"5F",X"13",X"05",X"16",X"64",X"5D",X"08",X"5E",X"A5",X"05",X"16",
		X"64",X"5D",X"08",X"5F",X"13",X"05",X"16",X"64",X"5D",X"08",X"5E",X"A5",X"05",X"16",X"64",X"5D",
		X"10",X"41",X"DB",X"05",X"10",X"63",X"F4",X"10",X"41",X"8B",X"05",X"10",X"64",X"5D",X"10",X"43",
		X"89",X"07",X"19",X"63",X"FE",X"10",X"3E",X"56",X"07",X"19",X"64",X"08",X"10",X"3F",X"05",X"07",
		X"19",X"64",X"5D",X"10",X"45",X"96",X"07",X"19",X"64",X"12",X"10",X"40",X"2D",X"07",X"19",X"64",
		X"1C",X"10",X"40",X"DC",X"07",X"19",X"64",X"5D",X"10",X"00",X"8D",X"06",X"10",X"64",X"68",X"10",
		X"00",X"2D",X"06",X"10",X"64",X"5D",X"10",X"00",X"8D",X"06",X"10",X"64",X"72",X"10",X"00",X"2D",
		X"06",X"10",X"64",X"5D",X"8E",X"B0",X"31",X"20",X"08",X"8E",X"B0",X"35",X"20",X"03",X"8E",X"B0",
		X"39",X"1F",X"20",X"AE",X"84",X"27",X"11",X"E1",X"88",X"32",X"27",X"05",X"AE",X"88",X"1A",X"20",
		X"F4",X"6F",X"88",X"1D",X"10",X"AF",X"88",X"14",X"86",X"01",X"39",X"F8",X"AD",X"F8",X"B5",X"F8",
		X"B5",X"F8",X"B5",X"F8",X"B5",X"F8",X"B5",X"F8",X"B5",X"F8",X"B5",X"F8",X"B5",X"F8",X"B5",X"F8",
		X"B5",X"F8",X"B5",X"F8",X"B5",X"F8",X"B5",X"F8",X"B5",X"F8",X"B5",X"F8",X"B5",X"F8",X"B5",X"F8",
		X"B5",X"F8",X"B5",X"F8",X"B5",X"F8",X"B5",X"F8",X"B5",X"F8",X"B5",X"F8",X"AD",X"F8",X"B5",X"65",
		X"44",X"65",X"49",X"65",X"4E",X"DC",X"06",X"27",X"4F",X"8D",X"53",X"9B",X"05",X"19",X"97",X"05",
		X"1F",X"98",X"99",X"04",X"19",X"97",X"04",X"24",X"07",X"86",X"00",X"99",X"03",X"19",X"97",X"03",
		X"DC",X"45",X"27",X"32",X"DC",X"01",X"93",X"06",X"2E",X"27",X"D3",X"45",X"DD",X"01",X"CC",X"00",
		X"00",X"DD",X"06",X"0C",X"00",X"8E",X"EC",X"7F",X"9F",X"21",X"8E",X"70",X"71",X"BD",X"6F",X"D3",
		X"8E",X"A9",X"27",X"86",X"01",X"BD",X"7E",X"EA",X"8E",X"A9",X"2D",X"86",X"01",X"BD",X"7E",X"EA",
		X"39",X"DD",X"01",X"CC",X"00",X"00",X"DD",X"06",X"39",X"8D",X"03",X"1E",X"89",X"39",X"8E",X"B3",
		X"4C",X"3A",X"3A",X"48",X"27",X"11",X"10",X"8E",X"B5",X"4C",X"EC",X"A6",X"AB",X"84",X"19",X"1E",
		X"89",X"A9",X"01",X"19",X"1E",X"89",X"39",X"EC",X"84",X"39",X"85",X"F0",X"26",X"0A",X"85",X"0F",
		X"26",X"12",X"C5",X"F0",X"26",X"14",X"20",X"1E",X"34",X"02",X"44",X"44",X"44",X"44",X"8A",X"30",
		X"A7",X"80",X"35",X"02",X"84",X"0F",X"8A",X"30",X"A7",X"80",X"34",X"04",X"54",X"54",X"54",X"54",
		X"CA",X"30",X"E7",X"80",X"35",X"04",X"C4",X"0F",X"CA",X"30",X"E7",X"80",X"39",X"0D",X"9C",X"26",
		X"FB",X"86",X"11",X"20",X"02",X"86",X"44",X"8E",X"BB",X"B9",X"7E",X"DF",X"05",X"0D",X"9C",X"26",
		X"EB",X"86",X"11",X"8E",X"BF",X"00",X"7E",X"DF",X"05",X"CC",X"0F",X"07",X"FD",X"C8",X"86",X"DC",
		X"0A",X"80",X"0F",X"FD",X"C8",X"84",X"CC",X"00",X"12",X"B7",X"C8",X"81",X"F7",X"C8",X"80",X"C6",
		X"06",X"96",X"03",X"26",X"0A",X"C6",X"04",X"96",X"04",X"26",X"04",X"C6",X"02",X"96",X"05",X"85",
		X"F0",X"26",X"06",X"5A",X"85",X"0F",X"26",X"01",X"5A",X"D7",X"12",X"86",X"22",X"8E",X"BF",X"00",
		X"7E",X"DF",X"05",X"EE",X"E4",X"37",X"36",X"ED",X"A1",X"AB",X"41",X"19",X"1E",X"89",X"A9",X"C4",
		X"19",X"1E",X"89",X"30",X"1F",X"26",X"F0",X"33",X"42",X"EF",X"E4",X"39",X"97",X"5B",X"0F",X"F0",
		X"81",X"01",X"27",X"06",X"81",X"04",X"27",X"02",X"03",X"F0",X"34",X"76",X"48",X"48",X"48",X"26",
		X"0E",X"8E",X"C0",X"00",X"31",X"89",X"00",X"BF",X"C6",X"45",X"BD",X"7F",X"26",X"20",X"35",X"CE",
		X"67",X"1A",X"33",X"C6",X"34",X"40",X"EE",X"C4",X"10",X"8E",X"C0",X"00",X"8E",X"01",X"C0",X"86",
		X"05",X"BD",X"DF",X"A0",X"EE",X"E4",X"EE",X"42",X"8E",X"10",X"10",X"10",X"8E",X"A6",X"D5",X"BD",
		X"DF",X"A0",X"EE",X"E4",X"EE",X"44",X"10",X"8E",X"A7",X"D5",X"BD",X"DF",X"A0",X"35",X"40",X"EC",
		X"46",X"FD",X"BA",X"1B",X"CC",X"FF",X"82",X"F7",X"CB",X"40",X"B7",X"CB",X"60",X"BD",X"67",X"B2",
		X"35",X"F6",X"75",X"00",X"78",X"00",X"7C",X"00",X"00",X"00",X"75",X"C0",X"79",X"00",X"7D",X"00",
		X"FF",X"FF",X"76",X"80",X"7A",X"00",X"7E",X"00",X"01",X"01",X"77",X"40",X"7B",X"00",X"7F",X"00",
		X"02",X"02",X"54",X"54",X"54",X"34",X"04",X"44",X"44",X"C6",X"20",X"3D",X"EB",X"E0",X"39",X"1F",
		X"30",X"8D",X"EF",X"8E",X"B5",X"9A",X"30",X"8B",X"B6",X"BA",X"1A",X"A7",X"84",X"39",X"81",X"F0",
		X"24",X"0D",X"81",X"90",X"24",X"0D",X"8D",X"DA",X"10",X"8E",X"B5",X"9A",X"A6",X"AB",X"39",X"86",
		X"3C",X"20",X"FB",X"86",X"3E",X"20",X"F7",X"B7",X"BA",X"1A",X"C6",X"08",X"CE",X"05",X"34",X"8D",
		X"20",X"CE",X"05",X"3C",X"8D",X"1B",X"CE",X"05",X"44",X"8D",X"16",X"39",X"B7",X"BA",X"1A",X"C6",
		X"07",X"CE",X"71",X"34",X"8D",X"0B",X"CE",X"71",X"3C",X"8D",X"06",X"CE",X"71",X"44",X"8D",X"01",
		X"39",X"34",X"04",X"34",X"04",X"BD",X"67",X"4F",X"33",X"C9",X"04",X"00",X"6A",X"E4",X"26",X"F5",
		X"35",X"86",X"8E",X"B5",X"9A",X"31",X"89",X"04",X"7F",X"5F",X"BD",X"7F",X"26",X"86",X"34",X"B7",
		X"BA",X"1A",X"C6",X"08",X"CE",X"01",X"A4",X"8D",X"D8",X"CE",X"01",X"AC",X"8D",X"D3",X"CE",X"01",
		X"B4",X"8D",X"CE",X"C6",X"07",X"CE",X"75",X"A4",X"8D",X"C7",X"CE",X"75",X"AC",X"8D",X"C2",X"CE",
		X"75",X"B4",X"8D",X"BD",X"86",X"14",X"B7",X"BA",X"1A",X"C6",X"07",X"CE",X"01",X"B4",X"BD",X"69",
		X"73",X"86",X"16",X"B7",X"BA",X"1A",X"CE",X"8D",X"B4",X"BD",X"69",X"73",X"86",X"1C",X"B7",X"BA",
		X"1A",X"C6",X"0E",X"CE",X"01",X"04",X"BD",X"69",X"73",X"86",X"1E",X"B7",X"BA",X"1A",X"CE",X"8D",
		X"04",X"BD",X"69",X"73",X"86",X"24",X"B7",X"BA",X"1A",X"C6",X"24",X"CE",X"01",X"EC",X"BD",X"67",
		X"A1",X"CE",X"01",X"F4",X"BD",X"67",X"A1",X"86",X"26",X"B7",X"BA",X"1A",X"CE",X"1D",X"9C",X"C6",
		X"03",X"BD",X"69",X"73",X"CE",X"19",X"9C",X"C6",X"02",X"BD",X"69",X"73",X"86",X"28",X"B7",X"BA",
		X"1A",X"CE",X"79",X"9C",X"BD",X"69",X"73",X"CE",X"75",X"9C",X"C6",X"03",X"BD",X"69",X"73",X"86",
		X"36",X"B7",X"BA",X"1A",X"CE",X"19",X"94",X"C6",X"02",X"BD",X"67",X"A1",X"CE",X"75",X"94",X"BD",
		X"67",X"A1",X"86",X"2C",X"B7",X"BA",X"1A",X"C6",X"0C",X"CE",X"31",X"34",X"BD",X"67",X"A1",X"CE",
		X"31",X"3C",X"BD",X"67",X"A1",X"86",X"2E",X"B7",X"BA",X"1A",X"C6",X"03",X"CE",X"25",X"34",X"BD",
		X"67",X"A1",X"CE",X"25",X"3C",X"BD",X"67",X"A1",X"C6",X"04",X"CE",X"61",X"34",X"BD",X"67",X"A1",
		X"CE",X"61",X"3C",X"BD",X"67",X"A1",X"86",X"18",X"B7",X"BA",X"1A",X"C6",X"08",X"CE",X"21",X"5C",
		X"BD",X"69",X"73",X"CE",X"25",X"5C",X"BD",X"69",X"73",X"86",X"1A",X"B7",X"BA",X"1A",X"C6",X"08",
		X"CE",X"69",X"5C",X"BD",X"69",X"73",X"CE",X"6D",X"5C",X"BD",X"69",X"73",X"CE",X"71",X"5C",X"BD",
		X"69",X"73",X"96",X"5B",X"81",X"02",X"27",X"18",X"86",X"20",X"B7",X"BA",X"1A",X"C6",X"04",X"CE",
		X"29",X"64",X"BD",X"69",X"73",X"86",X"22",X"B7",X"BA",X"1A",X"CE",X"69",X"64",X"BD",X"69",X"73",
		X"96",X"F0",X"26",X"22",X"86",X"2A",X"BD",X"67",X"77",X"C6",X"01",X"CE",X"01",X"44",X"BD",X"67",
		X"A1",X"86",X"30",X"B7",X"BA",X"1A",X"C6",X"02",X"CE",X"21",X"4C",X"BD",X"69",X"73",X"CE",X"25",
		X"4C",X"BD",X"69",X"73",X"20",X"1A",X"86",X"2E",X"BD",X"67",X"77",X"86",X"3A",X"B7",X"BA",X"1A",
		X"C6",X"08",X"CE",X"05",X"4C",X"BD",X"67",X"A1",X"C6",X"09",X"CE",X"01",X"54",X"BD",X"67",X"A1",
		X"96",X"F0",X"26",X"20",X"86",X"2A",X"BD",X"67",X"8C",X"C6",X"01",X"CE",X"8D",X"44",X"BD",X"67",
		X"A1",X"86",X"32",X"B7",X"BA",X"1A",X"C6",X"02",X"CE",X"71",X"4C",X"8D",X"36",X"CE",X"75",X"4C",
		X"8D",X"31",X"20",X"1A",X"86",X"2E",X"BD",X"67",X"8C",X"86",X"3A",X"B7",X"BA",X"1A",X"C6",X"07",
		X"CE",X"71",X"4C",X"BD",X"67",X"A1",X"C6",X"08",X"CE",X"71",X"54",X"BD",X"67",X"A1",X"96",X"E4",
		X"27",X"08",X"10",X"8E",X"69",X"C0",X"86",X"02",X"20",X"06",X"10",X"8E",X"69",X"96",X"86",X"0E",
		X"8D",X"10",X"39",X"34",X"04",X"34",X"04",X"BD",X"67",X"4F",X"33",X"48",X"6A",X"E4",X"26",X"F7",
		X"35",X"86",X"34",X"02",X"6A",X"E4",X"2D",X"0C",X"EE",X"A1",X"A6",X"A0",X"B7",X"BA",X"1A",X"BD",
		X"67",X"4F",X"20",X"F0",X"35",X"82",X"15",X"34",X"02",X"15",X"3C",X"02",X"29",X"34",X"04",X"29",
		X"3C",X"04",X"31",X"3C",X"10",X"5D",X"3C",X"12",X"6D",X"34",X"08",X"6D",X"3C",X"08",X"85",X"34",
		X"0A",X"85",X"3C",X"0A",X"11",X"AC",X"0C",X"11",X"B4",X"0C",X"7D",X"AC",X"0E",X"7D",X"B4",X"0E",
		X"49",X"34",X"06",X"49",X"3C",X"06",X"86",X"05",X"A7",X"C8",X"1F",X"CC",X"6D",X"F8",X"ED",X"C8",
		X"40",X"CC",X"00",X"00",X"A7",X"4E",X"A7",X"C8",X"1D",X"ED",X"C8",X"34",X"ED",X"C8",X"36",X"A7",
		X"C8",X"38",X"A7",X"C8",X"44",X"A7",X"C8",X"45",X"A7",X"C8",X"4A",X"A7",X"C8",X"43",X"A7",X"C8",
		X"4B",X"ED",X"C8",X"4C",X"A7",X"C8",X"4E",X"B6",X"AF",X"FB",X"A7",X"C8",X"3C",X"A7",X"C8",X"3B",
		X"8E",X"6A",X"1F",X"AF",X"C8",X"3E",X"8E",X"6A",X"0C",X"AF",X"4A",X"39",X"A6",X"4E",X"27",X"04",
		X"BD",X"30",X"7C",X"39",X"A6",X"C8",X"4E",X"27",X"03",X"7E",X"6D",X"CB",X"6E",X"D8",X"3E",X"A6",
		X"C8",X"4B",X"27",X"03",X"7E",X"6D",X"9C",X"8E",X"6A",X"8F",X"AF",X"C8",X"3E",X"EC",X"C8",X"14",
		X"ED",X"C8",X"5E",X"E1",X"C8",X"32",X"25",X"2F",X"22",X"33",X"10",X"8E",X"00",X"00",X"A1",X"C8",
		X"30",X"26",X"2E",X"A6",X"C8",X"1D",X"26",X"44",X"A6",X"C8",X"43",X"26",X"0B",X"96",X"D5",X"84",
		X"07",X"8B",X"01",X"A7",X"C8",X"43",X"20",X"34",X"6A",X"C8",X"43",X"26",X"1B",X"86",X"FF",X"A7",
		X"C8",X"1D",X"BD",X"39",X"13",X"20",X"11",X"10",X"BE",X"AF",X"F9",X"20",X"04",X"10",X"BE",X"AF",
		X"F7",X"A1",X"C8",X"30",X"25",X"07",X"22",X"0A",X"8E",X"00",X"00",X"20",X"08",X"BE",X"AF",X"F9",
		X"20",X"03",X"BE",X"AF",X"F7",X"10",X"AF",X"C8",X"36",X"AF",X"C8",X"34",X"7E",X"6D",X"9B",X"8E",
		X"6B",X"D4",X"AF",X"C8",X"3E",X"A6",X"C8",X"30",X"E6",X"C8",X"32",X"BD",X"67",X"5E",X"A7",X"C8",
		X"38",X"27",X"08",X"A7",X"C8",X"16",X"8E",X"6A",X"AE",X"AF",X"4A",X"7E",X"6D",X"9B",X"A6",X"C8",
		X"16",X"8E",X"6E",X"36",X"AE",X"86",X"A6",X"C8",X"30",X"E6",X"C8",X"32",X"6E",X"84",X"10",X"A3",
		X"C8",X"5E",X"27",X"08",X"20",X"23",X"10",X"A3",X"C8",X"5E",X"26",X"25",X"AE",X"C8",X"4C",X"27",
		X"0C",X"CC",X"00",X"00",X"A7",X"88",X"4B",X"A7",X"88",X"4E",X"ED",X"88",X"4C",X"BD",X"F9",X"16",
		X"39",X"C1",X"EC",X"25",X"5D",X"C6",X"EC",X"20",X"3F",X"C1",X"B1",X"22",X"55",X"C6",X"B1",X"20",
		X"27",X"C1",X"39",X"25",X"04",X"C6",X"39",X"20",X"2F",X"C1",X"37",X"22",X"45",X"C6",X"37",X"20",
		X"17",X"C1",X"38",X"22",X"3D",X"C6",X"38",X"20",X"0F",X"C1",X"97",X"22",X"35",X"C6",X"98",X"8E",
		X"00",X"00",X"AF",X"C8",X"34",X"BD",X"39",X"2F",X"E7",X"C8",X"32",X"EC",X"C8",X"36",X"2A",X"22",
		X"CC",X"00",X"00",X"ED",X"C8",X"36",X"20",X"1A",X"E7",X"C8",X"32",X"EC",X"C8",X"36",X"2F",X"12",
		X"20",X"EE",X"C1",X"68",X"25",X"0C",X"C6",X"68",X"20",X"EE",X"C1",X"48",X"25",X"04",X"C6",X"48",
		X"20",X"E6",X"CC",X"6A",X"0C",X"ED",X"4A",X"39",X"A7",X"C8",X"30",X"EC",X"C8",X"34",X"2A",X"F2",
		X"CC",X"00",X"00",X"ED",X"C8",X"34",X"20",X"EA",X"A7",X"C8",X"30",X"EC",X"C8",X"34",X"2F",X"E2",
		X"20",X"EE",X"81",X"23",X"22",X"DC",X"86",X"23",X"20",X"DE",X"81",X"70",X"25",X"D4",X"86",X"70",
		X"20",X"E6",X"81",X"1D",X"22",X"CC",X"86",X"1D",X"20",X"CE",X"81",X"76",X"25",X"C4",X"86",X"76",
		X"20",X"D6",X"81",X"25",X"22",X"BC",X"86",X"25",X"8D",X"3C",X"20",X"BC",X"81",X"6E",X"25",X"B2",
		X"86",X"6E",X"8D",X"32",X"20",X"C2",X"81",X"27",X"22",X"A8",X"86",X"27",X"8D",X"28",X"20",X"A8",
		X"81",X"6C",X"25",X"9E",X"86",X"6C",X"8D",X"1E",X"20",X"AE",X"C6",X"10",X"E7",X"C8",X"14",X"E6",
		X"C8",X"32",X"E7",X"C8",X"15",X"86",X"01",X"20",X"8F",X"C6",X"80",X"E7",X"C8",X"14",X"E6",X"C8",
		X"32",X"E7",X"C8",X"15",X"20",X"92",X"D6",X"38",X"27",X"09",X"EC",X"C8",X"14",X"A7",X"C8",X"30",
		X"E7",X"C8",X"32",X"39",X"8E",X"6C",X"3E",X"AF",X"C8",X"3E",X"EC",X"C8",X"36",X"2D",X"28",X"26",
		X"1C",X"EC",X"C8",X"34",X"26",X"2F",X"6C",X"C8",X"4A",X"A6",X"C8",X"4A",X"81",X"08",X"25",X"4B",
		X"A6",X"C8",X"43",X"26",X"46",X"BD",X"39",X"2F",X"6F",X"C8",X"4A",X"20",X"3E",X"E3",X"C8",X"32",
		X"A1",X"C8",X"5F",X"22",X"0A",X"20",X"0B",X"E3",X"C8",X"32",X"A1",X"C8",X"5F",X"24",X"03",X"A6",
		X"C8",X"5F",X"ED",X"C8",X"32",X"6F",X"C8",X"4A",X"EC",X"C8",X"34",X"2D",X"0C",X"27",X"1C",X"E3",
		X"C8",X"30",X"A1",X"C8",X"5E",X"22",X"0E",X"20",X"0F",X"E3",X"C8",X"30",X"A1",X"C8",X"5E",X"25",
		X"04",X"81",X"F0",X"25",X"03",X"A6",X"C8",X"5E",X"ED",X"C8",X"30",X"7E",X"6D",X"9B",X"8E",X"6D",
		X"07",X"AF",X"C8",X"3E",X"EC",X"C8",X"34",X"BD",X"6C",X"91",X"A6",X"C8",X"32",X"81",X"A0",X"22",
		X"08",X"81",X"58",X"22",X"07",X"86",X"04",X"20",X"05",X"4F",X"20",X"02",X"86",X"02",X"AE",X"C8",
		X"40",X"AE",X"86",X"AF",X"42",X"8E",X"6E",X"32",X"AE",X"86",X"AF",X"46",X"8D",X"05",X"6C",X"4F",
		X"7E",X"6D",X"9B",X"A6",X"46",X"44",X"40",X"AB",X"C8",X"30",X"A7",X"44",X"86",X"2A",X"E6",X"C8",
		X"31",X"2D",X"02",X"86",X"0A",X"A7",X"40",X"A6",X"47",X"44",X"40",X"AB",X"C8",X"32",X"A7",X"45",
		X"39",X"2D",X"40",X"2E",X"1A",X"86",X"FF",X"A7",X"C8",X"44",X"A6",X"C8",X"4B",X"26",X"0A",X"96",
		X"F4",X"26",X"06",X"CC",X"6D",X"F2",X"7E",X"6C",X"F5",X"CC",X"6D",X"F8",X"7E",X"6C",X"F5",X"A6",
		X"C8",X"44",X"27",X"0A",X"6F",X"C8",X"44",X"86",X"02",X"A7",X"C8",X"45",X"20",X"0E",X"A6",X"C8",
		X"45",X"8B",X"FE",X"2A",X"04",X"8D",X"32",X"86",X"06",X"A7",X"C8",X"45",X"8E",X"6D",X"FE",X"EC",
		X"86",X"20",X"22",X"A6",X"C8",X"44",X"27",X"0A",X"6F",X"C8",X"44",X"86",X"02",X"A7",X"C8",X"45",
		X"20",X"0E",X"A6",X"C8",X"45",X"8B",X"FE",X"2A",X"04",X"8D",X"0E",X"86",X"06",X"A7",X"C8",X"45",
		X"8E",X"6E",X"18",X"EC",X"86",X"ED",X"C8",X"40",X"39",X"8E",X"70",X"CD",X"03",X"E9",X"2D",X"03",
		X"8E",X"70",X"D1",X"BD",X"6F",X"D3",X"39",X"8E",X"6A",X"1F",X"AF",X"C8",X"3E",X"DC",X"D5",X"10",
		X"93",X"D9",X"25",X"21",X"AE",X"C8",X"4C",X"26",X"1C",X"BE",X"B0",X"09",X"27",X"09",X"8D",X"60",
		X"27",X"15",X"AE",X"88",X"1A",X"26",X"F7",X"BE",X"B0",X"0D",X"27",X"09",X"8D",X"52",X"27",X"07",
		X"AE",X"88",X"1A",X"26",X"F7",X"20",X"64",X"A6",X"0E",X"26",X"FA",X"A6",X"88",X"4E",X"27",X"19",
		X"96",X"D5",X"81",X"3C",X"22",X"EF",X"CC",X"00",X"00",X"A7",X"88",X"4E",X"10",X"AE",X"88",X"4C",
		X"ED",X"A8",X"4C",X"A7",X"A8",X"4B",X"A7",X"A8",X"4E",X"A6",X"C8",X"30",X"E6",X"C8",X"32",X"ED",
		X"88",X"14",X"ED",X"C8",X"14",X"AF",X"C8",X"4C",X"86",X"0C",X"A7",X"C8",X"43",X"86",X"FF",X"A7",
		X"88",X"1E",X"6F",X"88",X"1D",X"A7",X"88",X"4B",X"EF",X"88",X"4C",X"6F",X"88",X"2B",X"20",X"B5",
		X"A6",X"88",X"30",X"A0",X"C8",X"30",X"2A",X"01",X"40",X"81",X"08",X"22",X"0E",X"A6",X"88",X"32",
		X"A0",X"C8",X"32",X"2A",X"01",X"40",X"81",X"10",X"22",X"01",X"4F",X"39",X"8E",X"6A",X"1F",X"AF",
		X"C8",X"3E",X"8D",X"04",X"6C",X"4F",X"20",X"F3",X"96",X"D5",X"81",X"E8",X"25",X"04",X"96",X"D6",
		X"20",X"01",X"4F",X"BD",X"6C",X"91",X"AE",X"C8",X"4C",X"A6",X"88",X"42",X"AE",X"C8",X"40",X"AE",
		X"86",X"AF",X"42",X"8E",X"6E",X"32",X"AE",X"86",X"AF",X"46",X"39",X"6F",X"C8",X"4E",X"AE",X"C8",
		X"4C",X"A6",X"88",X"30",X"E6",X"88",X"34",X"2B",X"04",X"9B",X"ED",X"20",X"02",X"9B",X"EC",X"A7",
		X"C8",X"30",X"E6",X"88",X"32",X"CB",X"05",X"E7",X"C8",X"32",X"8D",X"BC",X"BD",X"6C",X"73",X"6C",
		X"4F",X"39",X"25",X"50",X"2D",X"14",X"2F",X"60",X"2A",X"58",X"28",X"0C",X"30",X"E0",X"6E",X"0C",
		X"6E",X"12",X"6E",X"0C",X"6E",X"06",X"2B",X"07",X"2D",X"A7",X"31",X"40",X"2B",X"B6",X"2E",X"3A",
		X"31",X"A0",X"2C",X"65",X"2E",X"CD",X"32",X"00",X"6E",X"26",X"6E",X"2C",X"6E",X"26",X"6E",X"20",
		X"25",X"FF",X"28",X"9F",X"2F",X"C0",X"26",X"AE",X"29",X"32",X"30",X"20",X"27",X"5D",X"29",X"C5",
		X"30",X"80",X"07",X"19",X"07",X"15",X"06",X"10",X"6A",X"F1",X"6A",X"F9",X"6B",X"01",X"6A",X"F9",
		X"6A",X"F1",X"6A",X"E9",X"6A",X"E9",X"6B",X"01",X"6B",X"01",X"6A",X"BE",X"6A",X"BE",X"6B",X"82",
		X"6B",X"8C",X"6A",X"C6",X"6A",X"C6",X"6B",X"96",X"6B",X"A0",X"6A",X"E1",X"6B",X"72",X"6B",X"7A",
		X"6A",X"F1",X"6B",X"01",X"6A",X"F9",X"6B",X"62",X"6B",X"6A",X"6A",X"E9",X"6B",X"09",X"6B",X"32",
		X"6B",X"3A",X"6B",X"AA",X"6B",X"B9",X"BD",X"27",X"F8",X"8E",X"6E",X"BF",X"20",X"06",X"BD",X"27",
		X"F8",X"8E",X"6E",X"C6",X"BD",X"33",X"01",X"86",X"FF",X"97",X"A9",X"97",X"DC",X"10",X"8E",X"6E",
		X"D8",X"86",X"11",X"34",X"02",X"BD",X"27",X"9B",X"31",X"24",X"6A",X"E4",X"26",X"F7",X"35",X"82",
		X"6A",X"4E",X"2A",X"1A",X"AE",X"4C",X"A6",X"80",X"27",X"09",X"A7",X"4E",X"EC",X"81",X"AF",X"4C",
		X"ED",X"D4",X"39",X"A6",X"4F",X"27",X"03",X"7E",X"27",X"D0",X"AE",X"48",X"AF",X"4C",X"39",X"AE",
		X"4A",X"CC",X"6F",X"99",X"20",X"04",X"AE",X"4A",X"EC",X"02",X"ED",X"48",X"ED",X"4C",X"EC",X"84",
		X"ED",X"40",X"CC",X"6E",X"A0",X"ED",X"42",X"39",X"BC",X"DF",X"6F",X"1C",X"BC",X"E3",X"6F",X"23",
		X"BD",X"13",X"6F",X"2A",X"BC",X"FF",X"6F",X"31",X"BC",X"E5",X"6F",X"38",X"BD",X"03",X"6F",X"3F",
		X"BC",X"FD",X"6F",X"4C",X"BD",X"07",X"6F",X"53",X"BD",X"27",X"6F",X"5A",X"BD",X"25",X"6F",X"61",
		X"BD",X"23",X"6F",X"68",X"BD",X"33",X"6F",X"6F",X"BD",X"47",X"6F",X"76",X"BD",X"43",X"6F",X"7D",
		X"BD",X"3D",X"6F",X"84",X"BD",X"3F",X"6F",X"8B",X"BD",X"45",X"6F",X"92",X"08",X"00",X"00",X"0A",
		X"FF",X"FA",X"00",X"02",X"00",X"00",X"0A",X"0F",X"DD",X"00",X"07",X"F9",X"FD",X"07",X"0F",X"F0",
		X"00",X"07",X"0F",X"F0",X"07",X"F9",X"FD",X"00",X"04",X"00",X"00",X"09",X"ED",X"FE",X"00",X"08",
		X"00",X"00",X"08",X"EC",X"AF",X"08",X"EC",X"CF",X"08",X"EC",X"EF",X"00",X"08",X"00",X"00",X"08",
		X"0E",X"F0",X"00",X"05",X"00",X"00",X"0D",X"ED",X"FE",X"00",X"04",X"0F",X"88",X"14",X"0F",X"F8",
		X"00",X"08",X"0F",X"88",X"10",X"0F",X"F8",X"00",X"0C",X"0F",X"88",X"0C",X"0F",X"F8",X"00",X"10",
		X"0F",X"88",X"08",X"0F",X"F8",X"00",X"06",X"FF",X"FF",X"07",X"F3",X"E0",X"00",X"0C",X"FF",X"FF",
		X"04",X"FE",X"F0",X"00",X"08",X"00",X"00",X"0D",X"E0",X"EF",X"00",X"0A",X"00",X"00",X"0B",X"0C",
		X"EF",X"00",X"0D",X"00",X"00",X"08",X"0F",X"FF",X"00",X"02",X"AF",X"E1",X"02",X"AF",X"F3",X"02",
		X"CF",X"F8",X"05",X"FF",X"FF",X"04",X"CF",X"F8",X"04",X"AF",X"F3",X"04",X"AF",X"F1",X"05",X"AF",
		X"D1",X"05",X"AF",X"C1",X"05",X"AF",X"B1",X"05",X"AF",X"A1",X"06",X"AF",X"81",X"07",X"8D",X"71",
		X"09",X"58",X"50",X"0A",X"36",X"40",X"0B",X"23",X"30",X"78",X"00",X"00",X"78",X"00",X"00",X"78",
		X"00",X"00",X"00",X"34",X"06",X"EC",X"84",X"D1",X"AE",X"25",X"0C",X"0F",X"99",X"8D",X"2D",X"D7",
		X"AE",X"EC",X"02",X"DD",X"AF",X"97",X"B2",X"35",X"86",X"96",X"B2",X"27",X"1A",X"0A",X"B2",X"26",
		X"16",X"0A",X"B0",X"27",X"09",X"96",X"AF",X"97",X"B2",X"96",X"B1",X"8D",X"0F",X"39",X"CC",X"00",
		X"FF",X"D7",X"99",X"97",X"AE",X"8D",X"05",X"39",X"0D",X"99",X"27",X"1B",X"97",X"B1",X"34",X"10",
		X"8E",X"70",X"E1",X"A6",X"86",X"B7",X"C9",X"82",X"B6",X"C9",X"83",X"84",X"F7",X"B7",X"C9",X"83",
		X"8A",X"08",X"B7",X"C9",X"83",X"35",X"90",X"39",X"34",X"06",X"CC",X"00",X"FF",X"7D",X"A9",X"04",
		X"27",X"0B",X"97",X"AE",X"D7",X"99",X"F4",X"A9",X"18",X"D7",X"9D",X"35",X"86",X"97",X"B2",X"97",
		X"99",X"97",X"9D",X"D7",X"AE",X"8D",X"C5",X"35",X"86",X"00",X"FF",X"0A",X"01",X"10",X"FF",X"5A",
		X"01",X"01",X"FF",X"14",X"01",X"04",X"FA",X"2D",X"01",X"61",X"F9",X"5A",X"01",X"1B",X"F8",X"FF",
		X"01",X"44",X"F8",X"3C",X"01",X"54",X"F8",X"78",X"01",X"0D",X"F0",X"B4",X"01",X"03",X"DC",X"10",
		X"03",X"06",X"CF",X"14",X"01",X"07",X"CF",X"14",X"01",X"1B",X"CD",X"3C",X"01",X"18",X"C8",X"5A",
		X"01",X"19",X"C8",X"5A",X"01",X"09",X"C3",X"46",X"01",X"30",X"BE",X"2D",X"01",X"01",X"BB",X"06",
		X"01",X"02",X"AA",X"0F",X"01",X"01",X"B4",X"06",X"01",X"40",X"B4",X"5A",X"01",X"43",X"B4",X"3C",
		X"01",X"12",X"AA",X"1E",X"01",X"1A",X"AA",X"2D",X"01",X"1F",X"A0",X"0F",X"01",X"62",X"9B",X"14",
		X"01",X"13",X"96",X"0A",X"01",X"14",X"96",X"0A",X"01",X"17",X"8C",X"0A",X"01",X"15",X"8C",X"14",
		X"01",X"60",X"8C",X"0A",X"01",X"16",X"82",X"78",X"01",X"1C",X"64",X"0A",X"01",X"1D",X"64",X"02",
		X"01",X"1E",X"64",X"02",X"01",X"08",X"3C",X"10",X"01",X"0B",X"0A",X"03",X"01",X"03",X"0A",X"3C",
		X"01",X"00",X"57",X"37",X"3E",X"08",X"05",X"21",X"10",X"1C",X"30",X"0A",X"23",X"0C",X"11",X"0E",
		X"0F",X"55",X"55",X"12",X"40",X"43",X"05",X"4C",X"37",X"2D",X"4E",X"17",X"53",X"3C",X"41",X"41",
		X"07",X"1F",X"14",X"27",X"52",X"08",X"25",X"26",X"28",X"28",X"29",X"2A",X"4D",X"25",X"25",X"2E",
		X"2F",X"39",X"31",X"32",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",
		X"00",X"3D",X"3D",X"3D",X"1C",X"0C",X"0C",X"0C",X"3D",X"33",X"49",X"4A",X"4B",X"4C",X"4D",X"4E",
		X"4F",X"50",X"51",X"52",X"53",X"0C",X"12",X"36",X"0A",X"00",X"00",X"01",X"02",X"04",X"08",X"10",
		X"20",X"3A",X"14",X"38",X"34",X"42",X"B6",X"B0",X"50",X"81",X"02",X"24",X"21",X"BD",X"F8",X"AD",
		X"26",X"1C",X"CC",X"02",X"00",X"ED",X"40",X"86",X"28",X"A7",X"4C",X"C6",X"04",X"86",X"02",X"ED",
		X"C8",X"46",X"6F",X"4D",X"AE",X"61",X"AF",X"C8",X"39",X"8E",X"71",X"70",X"AF",X"4A",X"35",X"C2",
		X"10",X"AE",X"C8",X"39",X"E6",X"A8",X"34",X"26",X"04",X"AD",X"D8",X"22",X"39",X"8E",X"70",X"D5",
		X"BD",X"6F",X"D3",X"8E",X"72",X"5D",X"A6",X"26",X"E6",X"86",X"EB",X"25",X"E7",X"45",X"A6",X"A8",
		X"34",X"2A",X"29",X"8E",X"A6",X"D5",X"3A",X"A6",X"84",X"A7",X"C8",X"44",X"A6",X"24",X"2B",X"D9",
		X"A1",X"C8",X"44",X"23",X"D4",X"8E",X"1A",X"B4",X"AF",X"C8",X"48",X"8E",X"1A",X"BD",X"AF",X"C8",
		X"4A",X"8E",X"1A",X"C6",X"AF",X"C8",X"4C",X"8E",X"71",X"FB",X"20",X"29",X"8E",X"A7",X"D5",X"3A",
		X"A6",X"84",X"80",X"09",X"A7",X"C8",X"44",X"A6",X"24",X"AB",X"26",X"A1",X"C8",X"44",X"24",X"A9",
		X"8E",X"1A",X"99",X"AF",X"C8",X"48",X"8E",X"1A",X"A2",X"AF",X"C8",X"4A",X"8E",X"1A",X"AB",X"AF",
		X"C8",X"4C",X"8E",X"72",X"0A",X"A7",X"44",X"5F",X"ED",X"C8",X"30",X"AF",X"4A",X"86",X"01",X"A7",
		X"C8",X"1F",X"CC",X"09",X"01",X"ED",X"46",X"BD",X"41",X"10",X"39",X"EC",X"C8",X"30",X"C3",X"FE",
		X"80",X"2B",X"2A",X"A1",X"C8",X"44",X"23",X"25",X"20",X"0B",X"EC",X"C8",X"30",X"C3",X"01",X"80",
		X"A1",X"C8",X"44",X"24",X"18",X"ED",X"C8",X"30",X"A7",X"44",X"A6",X"40",X"84",X"DF",X"6D",X"C8",
		X"31",X"2A",X"02",X"8A",X"20",X"A7",X"40",X"6C",X"4F",X"8D",X"09",X"27",X"03",X"AD",X"D8",X"22",
		X"BD",X"41",X"10",X"39",X"BE",X"B0",X"15",X"26",X"01",X"39",X"EC",X"04",X"E1",X"45",X"22",X"17",
		X"A1",X"44",X"22",X"13",X"E3",X"06",X"E1",X"45",X"25",X"0D",X"A1",X"44",X"25",X"09",X"A6",X"0E",
		X"26",X"05",X"6A",X"0E",X"8A",X"FF",X"39",X"AE",X"88",X"1A",X"26",X"DE",X"39",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"08",X"00",X"0A",X"00",X"00",X"00",X"CE",X"78",X"5B",
		X"10",X"8E",X"BB",X"A7",X"8E",X"00",X"10",X"BD",X"7F",X"33",X"39",X"86",X"01",X"A7",X"C8",X"1F",
		X"6F",X"C8",X"57",X"BD",X"63",X"23",X"AF",X"C8",X"54",X"6F",X"C8",X"56",X"11",X"A3",X"88",X"54",
		X"26",X"0A",X"A6",X"88",X"56",X"2B",X"02",X"86",X"01",X"A7",X"C8",X"56",X"CC",X"77",X"AF",X"ED",
		X"C8",X"40",X"CC",X"00",X"00",X"A7",X"4E",X"A7",X"C8",X"1D",X"A7",X"C8",X"2B",X"ED",X"C8",X"2C",
		X"ED",X"C8",X"34",X"ED",X"C8",X"36",X"ED",X"C8",X"47",X"A7",X"C8",X"38",X"A7",X"C8",X"3A",X"A7",
		X"C8",X"42",X"A7",X"C8",X"45",X"A7",X"C8",X"49",X"A7",X"C8",X"46",X"A7",X"C8",X"4A",X"A7",X"C8",
		X"4B",X"ED",X"C8",X"4C",X"A7",X"C8",X"4E",X"A7",X"C8",X"4F",X"B6",X"BB",X"B7",X"A7",X"C8",X"3C",
		X"A7",X"C8",X"3B",X"8E",X"73",X"09",X"AF",X"C8",X"3E",X"8E",X"72",X"EF",X"AF",X"4A",X"39",X"6E",
		X"D8",X"3E",X"A6",X"C8",X"2B",X"27",X"11",X"6A",X"C8",X"2B",X"26",X"0C",X"EC",X"C8",X"2C",X"ED",
		X"C8",X"14",X"6F",X"C8",X"1D",X"6F",X"C8",X"1E",X"39",X"A6",X"4E",X"27",X"28",X"AE",X"C8",X"4C",
		X"27",X"0C",X"CC",X"00",X"00",X"ED",X"88",X"4C",X"A7",X"88",X"4B",X"A7",X"88",X"4E",X"AE",X"C8",
		X"54",X"27",X"0E",X"A6",X"C8",X"56",X"27",X"09",X"CC",X"00",X"00",X"ED",X"88",X"54",X"A7",X"88",
		X"56",X"BD",X"30",X"7C",X"39",X"8E",X"74",X"2B",X"AF",X"C8",X"3E",X"8D",X"B5",X"FC",X"BB",X"9F",
		X"6D",X"C8",X"4E",X"27",X"03",X"CC",X"02",X"00",X"FD",X"BB",X"A3",X"CC",X"00",X"00",X"B3",X"BB",
		X"A3",X"FD",X"BB",X"A5",X"EC",X"C8",X"14",X"ED",X"C8",X"5E",X"0D",X"39",X"27",X"21",X"AE",X"C8",
		X"4C",X"27",X"12",X"CC",X"00",X"00",X"A7",X"C8",X"4E",X"ED",X"C8",X"4C",X"ED",X"88",X"4C",X"A7",
		X"88",X"4B",X"A7",X"88",X"4E",X"8E",X"00",X"00",X"10",X"8E",X"00",X"00",X"7E",X"74",X"21",X"E1",
		X"C8",X"32",X"25",X"3A",X"22",X"3E",X"10",X"8E",X"00",X"00",X"A1",X"C8",X"30",X"25",X"45",X"22",
		X"3E",X"A6",X"C8",X"1D",X"10",X"26",X"00",X"90",X"86",X"FF",X"A7",X"C8",X"1D",X"BD",X"39",X"13",
		X"A6",X"C8",X"4B",X"27",X"14",X"8E",X"70",X"A9",X"BD",X"6F",X"D3",X"AE",X"C8",X"4C",X"27",X"09",
		X"A7",X"88",X"4B",X"A7",X"C8",X"4E",X"6F",X"C8",X"4B",X"8E",X"00",X"00",X"20",X"19",X"10",X"BE",
		X"BB",X"A5",X"20",X"04",X"10",X"BE",X"BB",X"A3",X"A1",X"C8",X"30",X"25",X"07",X"27",X"EA",X"BE",
		X"BB",X"A3",X"20",X"03",X"BE",X"BB",X"A5",X"A6",X"C8",X"1D",X"26",X"45",X"E6",X"C8",X"49",X"26",
		X"05",X"8C",X"00",X"00",X"26",X"3B",X"EC",X"C8",X"36",X"27",X"0D",X"A6",X"C8",X"32",X"A0",X"C8",
		X"15",X"2A",X"01",X"40",X"81",X"04",X"22",X"05",X"6F",X"C8",X"49",X"20",X"24",X"86",X"FF",X"A7",
		X"C8",X"49",X"A6",X"C8",X"46",X"4A",X"2A",X"09",X"63",X"C8",X"3A",X"96",X"D5",X"84",X"03",X"8B",
		X"02",X"A7",X"C8",X"46",X"A6",X"C8",X"3A",X"2D",X"05",X"BE",X"BB",X"A3",X"20",X"03",X"BE",X"BB",
		X"A5",X"AF",X"C8",X"34",X"10",X"AF",X"C8",X"36",X"7E",X"77",X"AE",X"8E",X"76",X"5D",X"AF",X"C8",
		X"3E",X"A6",X"C8",X"30",X"E6",X"C8",X"32",X"BD",X"67",X"5E",X"A7",X"C8",X"38",X"27",X"08",X"A7",
		X"C8",X"16",X"8E",X"74",X"4A",X"AF",X"4A",X"7E",X"77",X"AE",X"A6",X"C8",X"16",X"8E",X"77",X"F3",
		X"AE",X"86",X"A6",X"C8",X"30",X"E6",X"C8",X"32",X"10",X"A3",X"C8",X"5E",X"26",X"09",X"6D",X"C8",
		X"56",X"2D",X"04",X"1A",X"04",X"6E",X"84",X"1C",X"FB",X"6E",X"84",X"10",X"26",X"01",X"13",X"CC",
		X"14",X"30",X"7E",X"74",X"CB",X"10",X"26",X"01",X"11",X"CC",X"26",X"30",X"20",X"4D",X"10",X"26",
		X"01",X"10",X"CC",X"46",X"30",X"20",X"44",X"10",X"26",X"00",X"FF",X"CC",X"6B",X"30",X"20",X"3B",
		X"10",X"26",X"00",X"EE",X"CC",X"83",X"30",X"20",X"32",X"10",X"26",X"00",X"DD",X"C6",X"A1",X"8E",
		X"78",X"6B",X"20",X"2E",X"10",X"26",X"00",X"D2",X"C6",X"A1",X"8E",X"78",X"83",X"20",X"23",X"10",
		X"26",X"00",X"DF",X"C6",X"31",X"8E",X"78",X"9B",X"20",X"18",X"10",X"26",X"00",X"D4",X"C6",X"31",
		X"8E",X"78",X"AB",X"20",X"0D",X"CC",X"72",X"EF",X"ED",X"4A",X"39",X"8E",X"BB",X"A7",X"A7",X"01",
		X"A7",X"09",X"E7",X"45",X"20",X"60",X"6A",X"C8",X"1C",X"26",X"70",X"8E",X"BB",X"AF",X"20",X"56",
		X"6A",X"C8",X"1C",X"26",X"66",X"8E",X"78",X"73",X"20",X"4C",X"6A",X"C8",X"1C",X"26",X"5C",X"8E",
		X"78",X"7B",X"20",X"42",X"6A",X"C8",X"1C",X"26",X"52",X"8E",X"78",X"8B",X"20",X"38",X"6A",X"C8",
		X"1C",X"26",X"48",X"8E",X"78",X"93",X"20",X"2E",X"10",X"26",X"01",X"07",X"0D",X"E4",X"10",X"26",
		X"01",X"01",X"8E",X"78",X"3B",X"20",X"1F",X"10",X"26",X"01",X"08",X"8E",X"78",X"4B",X"20",X"16",
		X"10",X"26",X"00",X"F7",X"0D",X"E4",X"10",X"26",X"00",X"F1",X"8E",X"78",X"33",X"20",X"07",X"10",
		X"26",X"00",X"F8",X"8E",X"78",X"43",X"EC",X"81",X"A7",X"C8",X"1C",X"E7",X"44",X"EC",X"81",X"ED",
		X"42",X"6C",X"4F",X"EC",X"81",X"ED",X"46",X"EC",X"84",X"ED",X"4A",X"39",X"6A",X"C8",X"1C",X"26",
		X"FA",X"8E",X"78",X"53",X"20",X"E0",X"6A",X"C8",X"1C",X"26",X"F0",X"8E",X"78",X"A3",X"20",X"D6",
		X"6A",X"C8",X"1C",X"26",X"E6",X"8E",X"78",X"B3",X"20",X"CC",X"27",X"E5",X"20",X"0C",X"27",X"E1",
		X"20",X"10",X"C1",X"EC",X"25",X"5D",X"C6",X"EC",X"20",X"3F",X"C1",X"B1",X"22",X"55",X"C6",X"B1",
		X"20",X"27",X"C1",X"39",X"25",X"04",X"C6",X"39",X"20",X"2F",X"C1",X"37",X"22",X"45",X"C6",X"37",
		X"20",X"17",X"C1",X"38",X"22",X"3D",X"C6",X"38",X"20",X"0F",X"C1",X"97",X"22",X"35",X"C6",X"98",
		X"8E",X"00",X"00",X"AF",X"C8",X"34",X"BD",X"39",X"2F",X"E7",X"C8",X"32",X"EC",X"C8",X"36",X"2A",
		X"22",X"CC",X"00",X"00",X"ED",X"C8",X"36",X"20",X"1A",X"E7",X"C8",X"32",X"EC",X"C8",X"36",X"2F",
		X"12",X"20",X"EE",X"C1",X"68",X"25",X"0C",X"C6",X"68",X"20",X"EE",X"C1",X"48",X"25",X"04",X"C6",
		X"48",X"20",X"E6",X"CC",X"72",X"EF",X"ED",X"4A",X"39",X"A7",X"C8",X"30",X"EC",X"C8",X"34",X"2A",
		X"F2",X"CC",X"00",X"00",X"ED",X"C8",X"34",X"20",X"EA",X"A7",X"C8",X"30",X"EC",X"C8",X"34",X"2F",
		X"E2",X"20",X"EE",X"81",X"24",X"22",X"DC",X"86",X"24",X"20",X"DE",X"81",X"70",X"25",X"D4",X"86",
		X"70",X"20",X"E6",X"81",X"1E",X"22",X"CC",X"86",X"1E",X"20",X"CE",X"81",X"74",X"25",X"C4",X"86",
		X"74",X"20",X"D6",X"81",X"27",X"22",X"BC",X"86",X"27",X"20",X"BE",X"81",X"6C",X"25",X"B4",X"86",
		X"6C",X"20",X"C6",X"81",X"28",X"22",X"AC",X"86",X"28",X"20",X"AE",X"81",X"6C",X"25",X"A4",X"86",
		X"6C",X"20",X"B6",X"C6",X"10",X"E7",X"C8",X"14",X"E6",X"C8",X"32",X"E7",X"C8",X"15",X"C6",X"FF",
		X"E7",X"C8",X"1E",X"86",X"01",X"20",X"92",X"C6",X"80",X"E7",X"C8",X"14",X"E6",X"C8",X"32",X"E7",
		X"C8",X"15",X"C6",X"FF",X"E7",X"C8",X"1E",X"20",X"90",X"BD",X"38",X"52",X"39",X"8E",X"76",X"ED",
		X"AF",X"C8",X"3E",X"A6",X"C8",X"4E",X"27",X"06",X"AE",X"C8",X"4C",X"A7",X"88",X"4E",X"A6",X"C8",
		X"48",X"BB",X"BB",X"B8",X"A7",X"C8",X"48",X"24",X"0B",X"6C",X"C8",X"47",X"6A",X"C8",X"3C",X"2A",
		X"03",X"6F",X"C8",X"3C",X"EC",X"C8",X"36",X"2D",X"20",X"26",X"14",X"EC",X"C8",X"34",X"26",X"27",
		X"6C",X"C8",X"4A",X"A6",X"C8",X"4A",X"81",X"08",X"25",X"20",X"BD",X"39",X"2F",X"20",X"18",X"E3",
		X"C8",X"32",X"A1",X"C8",X"5F",X"22",X"0A",X"20",X"0B",X"E3",X"C8",X"32",X"A1",X"C8",X"5F",X"24",
		X"03",X"A6",X"C8",X"5F",X"ED",X"C8",X"32",X"6F",X"C8",X"4A",X"A6",X"C8",X"49",X"27",X"08",X"EC",
		X"C8",X"34",X"E3",X"C8",X"30",X"20",X"20",X"EC",X"C8",X"34",X"2D",X"0C",X"27",X"1C",X"E3",X"C8",
		X"30",X"A1",X"C8",X"5E",X"22",X"0E",X"20",X"0F",X"E3",X"C8",X"30",X"A1",X"C8",X"5E",X"25",X"04",
		X"81",X"F0",X"25",X"03",X"A6",X"C8",X"5E",X"ED",X"C8",X"30",X"7E",X"77",X"AE",X"8E",X"77",X"A0",
		X"AF",X"C8",X"3E",X"96",X"39",X"27",X"05",X"CC",X"77",X"AF",X"20",X"37",X"EC",X"C8",X"34",X"2D",
		X"22",X"2E",X"13",X"96",X"D5",X"2D",X"24",X"20",X"15",X"A6",X"C8",X"45",X"8B",X"FE",X"2A",X"02",
		X"86",X"06",X"A7",X"C8",X"45",X"39",X"8D",X"F1",X"96",X"D6",X"81",X"E0",X"22",X"0D",X"8E",X"77",
		X"B5",X"20",X"0B",X"8D",X"E4",X"96",X"D6",X"81",X"E0",X"22",X"F3",X"8E",X"77",X"CF",X"A6",X"C8",
		X"45",X"EC",X"86",X"ED",X"C8",X"40",X"A6",X"C8",X"32",X"81",X"A0",X"22",X"09",X"81",X"58",X"22",
		X"0A",X"CC",X"04",X"06",X"20",X"08",X"CC",X"00",X"00",X"20",X"03",X"CC",X"02",X"00",X"A7",X"C8",
		X"42",X"E7",X"C8",X"2A",X"8E",X"77",X"E9",X"AE",X"86",X"AF",X"46",X"AE",X"C8",X"40",X"AE",X"86",
		X"AF",X"42",X"8E",X"77",X"EF",X"30",X"86",X"DC",X"D5",X"10",X"A3",X"84",X"25",X"03",X"BD",X"71",
		X"44",X"A6",X"46",X"44",X"40",X"AB",X"C8",X"30",X"A7",X"44",X"86",X"2A",X"E6",X"C8",X"31",X"2D",
		X"02",X"86",X"0A",X"A7",X"40",X"A6",X"47",X"44",X"40",X"AB",X"C8",X"32",X"A7",X"45",X"6C",X"4F",
		X"A6",X"C8",X"56",X"2A",X"19",X"AE",X"C8",X"54",X"A6",X"C8",X"42",X"A7",X"88",X"3B",X"20",X"0E",
		X"6A",X"C8",X"3B",X"2A",X"09",X"A6",X"C8",X"3C",X"A7",X"C8",X"3B",X"7E",X"73",X"09",X"39",X"63",
		X"05",X"6A",X"2B",X"6F",X"59",X"77",X"C3",X"77",X"C9",X"77",X"C3",X"77",X"BD",X"64",X"31",X"6A",
		X"FD",X"6F",X"FB",X"65",X"5D",X"6B",X"CF",X"70",X"9D",X"66",X"89",X"6C",X"A1",X"71",X"3F",X"77",
		X"DD",X"77",X"E3",X"77",X"DD",X"77",X"D7",X"5F",X"81",X"67",X"B5",X"6D",X"73",X"60",X"AD",X"68",
		X"87",X"6E",X"15",X"61",X"D9",X"69",X"59",X"6E",X"B7",X"0C",X"19",X"0A",X"15",X"09",X"12",X"FC",
		X"00",X"F8",X"00",X"FD",X"80",X"74",X"6B",X"74",X"75",X"74",X"7E",X"74",X"87",X"74",X"90",X"74",
		X"99",X"74",X"A4",X"74",X"AF",X"74",X"BA",X"75",X"6A",X"75",X"6A",X"75",X"08",X"75",X"20",X"75",
		X"6E",X"75",X"6E",X"75",X"17",X"75",X"2F",X"75",X"72",X"76",X"03",X"76",X"0B",X"75",X"82",X"75",
		X"92",X"75",X"8A",X"75",X"F3",X"75",X"FB",X"75",X"7A",X"75",X"9A",X"75",X"C3",X"75",X"CB",X"76",
		X"33",X"76",X"47",X"08",X"6C",X"5F",X"13",X"05",X"16",X"75",X"4C",X"08",X"21",X"5E",X"A5",X"05",
		X"16",X"75",X"4C",X"08",X"6B",X"5F",X"13",X"05",X"16",X"75",X"4C",X"08",X"23",X"5E",X"A5",X"05",
		X"16",X"75",X"4C",X"14",X"21",X"5F",X"81",X"01",X"01",X"76",X"59",X"10",X"00",X"41",X"8B",X"05",
		X"10",X"74",X"D6",X"10",X"00",X"41",X"DB",X"05",X"10",X"75",X"4C",X"10",X"10",X"42",X"2B",X"07",
		X"19",X"74",X"E0",X"10",X"10",X"42",X"DA",X"07",X"19",X"74",X"EA",X"10",X"10",X"43",X"89",X"07",
		X"19",X"75",X"4C",X"10",X"7D",X"44",X"38",X"07",X"19",X"74",X"F4",X"10",X"7D",X"44",X"E7",X"07",
		X"19",X"74",X"FE",X"10",X"7D",X"45",X"96",X"07",X"19",X"75",X"4C",X"10",X"31",X"00",X"2D",X"06",
		X"10",X"75",X"56",X"10",X"32",X"00",X"8D",X"06",X"10",X"75",X"4C",X"10",X"5C",X"00",X"2D",X"06",
		X"10",X"75",X"60",X"10",X"5B",X"00",X"8D",X"06",X"10",X"75",X"4C",X"1A",X"50",X"BD",X"E0",X"EC",
		X"C6",X"0A",X"BD",X"E5",X"61",X"1C",X"AF",X"BD",X"DB",X"41",X"0F",X"60",X"8E",X"79",X"60",X"BD",
		X"F5",X"42",X"8E",X"79",X"66",X"BD",X"F5",X"4F",X"CC",X"33",X"0E",X"B7",X"BC",X"CD",X"B7",X"BC",
		X"D4",X"F7",X"BC",X"CE",X"8E",X"00",X"26",X"BF",X"BC",X"CA",X"C6",X"35",X"F7",X"BC",X"CC",X"F7",
		X"BC",X"D3",X"CE",X"79",X"6C",X"AE",X"C1",X"BF",X"BC",X"C8",X"8E",X"BC",X"C8",X"BD",X"F5",X"42",
		X"10",X"AE",X"C1",X"8E",X"00",X"DA",X"A6",X"C4",X"30",X"86",X"BF",X"BC",X"D1",X"8E",X"BC",X"D5",
		X"BF",X"BC",X"CF",X"A6",X"22",X"BD",X"4B",X"4E",X"A6",X"21",X"BD",X"4B",X"51",X"A6",X"C0",X"27",
		X"07",X"7C",X"A6",X"4B",X"86",X"3A",X"A7",X"80",X"A6",X"A4",X"BD",X"4B",X"51",X"A6",X"1F",X"81",
		X"20",X"26",X"04",X"86",X"30",X"A7",X"1F",X"86",X"FF",X"A7",X"84",X"8E",X"BC",X"CF",X"BD",X"F5",
		X"42",X"F6",X"BC",X"CC",X"FB",X"BC",X"CE",X"F7",X"BC",X"CC",X"F7",X"BC",X"D3",X"AE",X"C1",X"26",
		X"A6",X"86",X"04",X"BD",X"E0",X"76",X"BD",X"E5",X"1F",X"96",X"60",X"27",X"F9",X"0F",X"60",X"39",
		X"79",X"A5",X"00",X"5C",X"21",X"11",X"79",X"B8",X"00",X"68",X"DF",X"22",X"79",X"CE",X"A9",X"1B",
		X"00",X"79",X"DE",X"A9",X"1E",X"00",X"79",X"F0",X"A9",X"21",X"00",X"7A",X"01",X"A9",X"24",X"00",
		X"7A",X"0E",X"A9",X"27",X"00",X"7A",X"24",X"A9",X"2A",X"FA",X"7A",X"3F",X"A9",X"2D",X"00",X"7A",
		X"50",X"A9",X"30",X"00",X"7A",X"64",X"A9",X"33",X"00",X"7A",X"75",X"A9",X"36",X"00",X"7A",X"8A",
		X"A9",X"39",X"FA",X"00",X"00",X"42",X"4F",X"4F",X"4B",X"4B",X"45",X"45",X"50",X"49",X"4E",X"47",
		X"20",X"54",X"4F",X"54",X"41",X"4C",X"53",X"FF",X"50",X"52",X"45",X"53",X"53",X"20",X"41",X"44",
		X"56",X"41",X"4E",X"43",X"45",X"20",X"54",X"4F",X"20",X"45",X"58",X"49",X"54",X"FF",X"4C",X"45",
		X"46",X"54",X"20",X"53",X"4C",X"4F",X"54",X"20",X"43",X"4F",X"49",X"4E",X"53",X"FF",X"43",X"45",
		X"4E",X"54",X"45",X"52",X"20",X"53",X"4C",X"4F",X"54",X"20",X"43",X"4F",X"49",X"4E",X"53",X"FF",
		X"52",X"49",X"47",X"48",X"54",X"20",X"53",X"4C",X"4F",X"54",X"20",X"43",X"4F",X"49",X"4E",X"53",
		X"FF",X"50",X"41",X"49",X"44",X"20",X"43",X"52",X"45",X"44",X"49",X"54",X"53",X"FF",X"45",X"58",
		X"54",X"52",X"41",X"20",X"4D",X"49",X"53",X"53",X"49",X"4F",X"4E",X"53",X"20",X"45",X"41",X"52",
		X"4E",X"45",X"44",X"FF",X"54",X"4F",X"54",X"41",X"4C",X"20",X"50",X"4C",X"41",X"59",X"20",X"54",
		X"49",X"4D",X"45",X"20",X"28",X"48",X"4F",X"55",X"52",X"3A",X"4D",X"49",X"4E",X"29",X"FF",X"54",
		X"4F",X"54",X"41",X"4C",X"20",X"4D",X"45",X"4E",X"20",X"50",X"4C",X"41",X"59",X"45",X"44",X"FF",
		X"54",X"4F",X"54",X"41",X"4C",X"20",X"53",X"49",X"4E",X"47",X"4C",X"45",X"20",X"50",X"4C",X"41",
		X"59",X"45",X"52",X"FF",X"54",X"4F",X"54",X"41",X"4C",X"20",X"54",X"57",X"4F",X"20",X"50",X"4C",
		X"41",X"59",X"45",X"52",X"FF",X"54",X"4F",X"54",X"41",X"4C",X"20",X"43",X"52",X"45",X"44",X"49",
		X"54",X"53",X"20",X"50",X"4C",X"41",X"59",X"45",X"44",X"FF",X"41",X"56",X"45",X"52",X"41",X"47",
		X"45",X"20",X"54",X"49",X"4D",X"45",X"2F",X"47",X"41",X"4D",X"45",X"20",X"28",X"4D",X"49",X"4E",
		X"3A",X"53",X"45",X"43",X"29",X"FF",X"86",X"4B",X"97",X"9A",X"8E",X"70",X"69",X"BD",X"6F",X"D3",
		X"96",X"E4",X"26",X"03",X"BD",X"00",X"B5",X"BD",X"E2",X"29",X"7F",X"A6",X"83",X"BD",X"6E",X"7E",
		X"10",X"8E",X"7D",X"B6",X"0F",X"39",X"BD",X"7C",X"25",X"BD",X"7C",X"AE",X"96",X"11",X"81",X"64",
		X"26",X"33",X"DC",X"45",X"FD",X"A6",X"84",X"4F",X"5F",X"DD",X"45",X"BD",X"3A",X"E6",X"34",X"01",
		X"1A",X"50",X"86",X"14",X"8E",X"7B",X"1A",X"BD",X"F8",X"FE",X"86",X"14",X"8E",X"7B",X"6A",X"BD",
		X"F8",X"FE",X"35",X"01",X"86",X"FF",X"97",X"9A",X"BD",X"7C",X"52",X"BD",X"29",X"1E",X"FC",X"A6",
		X"84",X"DD",X"45",X"20",X"06",X"BD",X"3A",X"71",X"BD",X"E5",X"1F",X"BD",X"7C",X"52",X"BD",X"27",
		X"7E",X"BD",X"33",X"01",X"BD",X"E5",X"1F",X"0F",X"9A",X"39",X"6F",X"45",X"CC",X"FF",X"FF",X"A7",
		X"4D",X"E7",X"C8",X"42",X"A7",X"C8",X"43",X"8E",X"7B",X"2D",X"AF",X"4A",X"39",X"6A",X"C8",X"43",
		X"26",X"0B",X"8E",X"70",X"5D",X"BD",X"6F",X"D3",X"86",X"08",X"A7",X"C8",X"43",X"6A",X"4D",X"26",
		X"20",X"86",X"02",X"A7",X"4D",X"CC",X"01",X"88",X"D3",X"06",X"DD",X"06",X"6A",X"C8",X"42",X"26",
		X"10",X"CC",X"00",X"28",X"D3",X"06",X"DD",X"06",X"86",X"C8",X"A7",X"4D",X"8E",X"7B",X"62",X"AF",
		X"4A",X"39",X"6A",X"4D",X"26",X"03",X"AD",X"D8",X"22",X"39",X"6F",X"45",X"CC",X"5A",X"12",X"A7",
		X"4D",X"E7",X"C8",X"42",X"8E",X"7B",X"7A",X"AF",X"4A",X"39",X"6A",X"4D",X"26",X"0F",X"86",X"2D",
		X"A7",X"4D",X"BD",X"00",X"B5",X"6A",X"C8",X"42",X"26",X"03",X"AD",X"D8",X"22",X"39",X"86",X"4B",
		X"97",X"9A",X"BD",X"E2",X"29",X"7F",X"A6",X"83",X"86",X"FF",X"97",X"DC",X"10",X"8E",X"7D",X"4A",
		X"0F",X"39",X"BD",X"7C",X"25",X"86",X"73",X"BD",X"E5",X"1F",X"4A",X"26",X"FA",X"73",X"A6",X"83",
		X"10",X"8E",X"7D",X"80",X"8D",X"6F",X"BD",X"E5",X"1F",X"BD",X"6E",X"76",X"BD",X"7C",X"AE",X"BD",
		X"3A",X"31",X"CC",X"00",X"3C",X"BD",X"3A",X"ED",X"BD",X"7C",X"52",X"BD",X"27",X"90",X"0F",X"9A",
		X"39",X"96",X"40",X"27",X"0D",X"96",X"2C",X"27",X"08",X"B6",X"BB",X"B9",X"27",X"03",X"BD",X"7E",
		X"73",X"39",X"DC",X"10",X"C3",X"00",X"01",X"DD",X"10",X"39",X"96",X"40",X"27",X"15",X"96",X"2C",
		X"27",X"11",X"96",X"09",X"48",X"8E",X"7C",X"04",X"AE",X"86",X"BD",X"F5",X"CC",X"CC",X"00",X"73",
		X"BD",X"3A",X"ED",X"39",X"3C",X"BA",X"3C",X"D0",X"96",X"40",X"27",X"0E",X"B6",X"A9",X"02",X"81",
		X"01",X"27",X"07",X"0A",X"00",X"CC",X"EC",X"77",X"DD",X"21",X"CC",X"EC",X"D5",X"DD",X"1D",X"CC",
		X"EC",X"FA",X"DD",X"1F",X"39",X"34",X"01",X"1A",X"50",X"BD",X"39",X"5D",X"BD",X"F9",X"F6",X"CC",
		X"00",X"00",X"DD",X"D5",X"86",X"FF",X"97",X"96",X"CE",X"90",X"00",X"BD",X"7C",X"90",X"CE",X"90",
		X"60",X"BD",X"7C",X"90",X"35",X"01",X"A6",X"9F",X"BB",X"1D",X"27",X"05",X"BD",X"E5",X"1F",X"20",
		X"F5",X"39",X"BD",X"E5",X"1F",X"8D",X"03",X"26",X"F9",X"39",X"BD",X"34",X"74",X"1A",X"50",X"CE",
		X"90",X"00",X"8D",X"44",X"CE",X"90",X"60",X"8D",X"3F",X"1C",X"AF",X"96",X"66",X"8E",X"B0",X"00",
		X"A0",X"88",X"54",X"A0",X"88",X"58",X"A0",X"88",X"60",X"A0",X"88",X"5C",X"39",X"6F",X"C8",X"27",
		X"7D",X"A6",X"83",X"27",X"07",X"AE",X"C8",X"28",X"27",X"02",X"AF",X"4A",X"A6",X"4C",X"AD",X"B6",
		X"EE",X"C8",X"12",X"26",X"E8",X"39",X"A6",X"4E",X"26",X"0E",X"A6",X"C8",X"30",X"81",X"01",X"23",
		X"04",X"81",X"8F",X"25",X"03",X"BD",X"F9",X"4B",X"EE",X"C8",X"12",X"26",X"E9",X"39",X"BD",X"E5",
		X"1F",X"BD",X"7C",X"5A",X"1A",X"50",X"CE",X"90",X"00",X"8D",X"19",X"26",X"05",X"CE",X"90",X"60",
		X"8D",X"12",X"1C",X"AF",X"26",X"E8",X"39",X"A6",X"45",X"81",X"AC",X"24",X"07",X"AB",X"47",X"81",
		X"60",X"23",X"01",X"39",X"EE",X"C8",X"12",X"26",X"EE",X"39",X"A6",X"4E",X"26",X"2E",X"8E",X"7D",
		X"0D",X"A6",X"C8",X"32",X"2B",X"05",X"5F",X"81",X"46",X"20",X"04",X"C6",X"01",X"81",X"B3",X"59",
		X"A6",X"C8",X"30",X"81",X"49",X"22",X"05",X"59",X"81",X"23",X"20",X"03",X"59",X"81",X"6E",X"59",
		X"58",X"AE",X"95",X"AF",X"C8",X"14",X"6F",X"C8",X"3C",X"6F",X"C8",X"1D",X"39",X"51",X"33",X"51",
		X"33",X"51",X"31",X"51",X"31",X"51",X"33",X"51",X"33",X"51",X"31",X"51",X"31",X"51",X"2B",X"51",
		X"2B",X"51",X"29",X"51",X"29",X"51",X"2B",X"51",X"2B",X"51",X"29",X"51",X"29",X"A6",X"4E",X"26",
		X"02",X"6C",X"4E",X"39",X"A6",X"4E",X"26",X"0B",X"AE",X"4A",X"AF",X"C8",X"28",X"8E",X"7D",X"EC",
		X"AF",X"4A",X"39",X"8E",X"00",X"00",X"AF",X"C8",X"28",X"39",X"7D",X"34",X"7D",X"34",X"7D",X"34",
		X"7D",X"34",X"7D",X"34",X"7D",X"34",X"7D",X"34",X"7D",X"34",X"7D",X"34",X"7D",X"34",X"7D",X"34",
		X"7D",X"38",X"7D",X"38",X"7D",X"38",X"7D",X"38",X"7D",X"38",X"7D",X"34",X"7D",X"34",X"7D",X"34",
		X"7D",X"38",X"7D",X"38",X"7D",X"34",X"7D",X"34",X"7D",X"34",X"7D",X"34",X"7D",X"34",X"7D",X"34",
		X"F9",X"4B",X"28",X"1B",X"28",X"1B",X"28",X"1B",X"28",X"1B",X"28",X"1B",X"28",X"1B",X"28",X"1B",
		X"28",X"1B",X"28",X"1B",X"7D",X"EC",X"28",X"1B",X"26",X"08",X"26",X"08",X"26",X"08",X"43",X"8C",
		X"28",X"1B",X"41",X"BB",X"7D",X"EC",X"28",X"1B",X"28",X"1B",X"49",X"9D",X"3D",X"D4",X"28",X"1B",
		X"7D",X"ED",X"F9",X"4B",X"F9",X"4B",X"F9",X"4B",X"7D",X"EC",X"7C",X"DA",X"7C",X"DA",X"7D",X"2D",
		X"7C",X"DA",X"7C",X"DA",X"7C",X"DA",X"7C",X"DA",X"28",X"1B",X"7D",X"EC",X"28",X"1B",X"26",X"08",
		X"26",X"08",X"26",X"08",X"43",X"8C",X"28",X"1B",X"41",X"BB",X"7D",X"EC",X"7D",X"EC",X"7D",X"EC",
		X"49",X"9D",X"3D",X"D4",X"28",X"1B",X"7D",X"ED",X"F9",X"4B",X"F9",X"4B",X"39",X"6D",X"4E",X"26",
		X"03",X"BD",X"28",X"1B",X"39",X"E6",X"2C",X"8E",X"B0",X"00",X"58",X"3A",X"6C",X"84",X"A6",X"03",
		X"27",X"02",X"0C",X"65",X"0C",X"66",X"CC",X"00",X"00",X"ED",X"A8",X"18",X"EE",X"01",X"EF",X"A8",
		X"1A",X"27",X"04",X"10",X"AF",X"C8",X"18",X"10",X"AF",X"01",X"39",X"34",X"40",X"E6",X"4C",X"8E",
		X"B0",X"00",X"58",X"3A",X"A6",X"03",X"27",X"02",X"0A",X"65",X"0A",X"66",X"6A",X"00",X"26",X"07",
		X"CC",X"00",X"00",X"ED",X"01",X"35",X"C0",X"10",X"AE",X"C8",X"18",X"26",X"0B",X"EE",X"C8",X"1A",
		X"EF",X"01",X"10",X"AF",X"C8",X"18",X"35",X"C0",X"AE",X"C8",X"1A",X"AF",X"A8",X"1A",X"27",X"04",
		X"10",X"AF",X"88",X"18",X"35",X"C0",X"C6",X"6C",X"8E",X"B0",X"00",X"6F",X"80",X"5A",X"26",X"FB",
		X"0F",X"65",X"0F",X"66",X"C6",X"FF",X"F7",X"B0",X"0B",X"F7",X"B0",X"0F",X"F7",X"B0",X"07",X"F7",
		X"B0",X"23",X"39",X"34",X"77",X"1A",X"50",X"8E",X"BF",X"00",X"10",X"8E",X"BB",X"B9",X"86",X"14",
		X"34",X"02",X"EC",X"84",X"EE",X"A4",X"ED",X"A1",X"EF",X"81",X"6A",X"E4",X"26",X"F4",X"35",X"02",
		X"35",X"F7",X"91",X"09",X"27",X"02",X"8D",X"DB",X"39",X"86",X"FF",X"B7",X"BC",X"2D",X"BD",X"DF",
		X"81",X"BD",X"ED",X"1E",X"BD",X"DE",X"03",X"CE",X"7F",X"69",X"8D",X"17",X"96",X"2C",X"26",X"0B",
		X"0F",X"00",X"CC",X"EC",X"F9",X"DD",X"21",X"DD",X"1D",X"DD",X"1F",X"8D",X"B6",X"CE",X"7F",X"42",
		X"8D",X"01",X"39",X"10",X"8E",X"BF",X"00",X"8E",X"00",X"27",X"8D",X"67",X"B6",X"A9",X"02",X"97",
		X"00",X"DC",X"45",X"DD",X"01",X"39",X"0A",X"0F",X"2A",X"0F",X"86",X"3B",X"97",X"0F",X"DC",X"0D",
		X"C3",X"00",X"01",X"DD",X"0D",X"24",X"02",X"0C",X"0C",X"39",X"AB",X"84",X"19",X"A7",X"80",X"24",
		X"10",X"86",X"00",X"A9",X"84",X"19",X"A7",X"80",X"24",X"07",X"86",X"00",X"A9",X"84",X"19",X"A7",
		X"84",X"39",X"34",X"02",X"AB",X"02",X"A7",X"02",X"A6",X"01",X"89",X"00",X"A7",X"01",X"A6",X"84",
		X"89",X"00",X"A7",X"84",X"35",X"82",X"34",X"06",X"EC",X"01",X"E3",X"21",X"ED",X"01",X"A6",X"84",
		X"A9",X"A4",X"A7",X"84",X"35",X"86",X"34",X"35",X"BD",X"DF",X"C4",X"E7",X"80",X"AC",X"64",X"23",
		X"F7",X"35",X"B5",X"34",X"75",X"BD",X"DF",X"C4",X"E6",X"C0",X"E7",X"A0",X"30",X"1F",X"26",X"F5",
		X"35",X"F5",X"00",X"27",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"96",X"00",X"00",
		X"00",X"3C",X"00",X"01",X"00",X"1D",X"9A",X"1D",X"7D",X"00",X"00",X"1D",X"83",X"00",X"00",X"EC",
		X"D5",X"EC",X"FA",X"EC",X"7F",X"A6",X"6A",X"00",X"00",X"00",X"27",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"8B",X"96",X"00",X"00",X"00",X"3C",X"00",X"01",X"00",X"72",X"9A",X"72",X"7D",
		X"00",X"00",X"72",X"83",X"00",X"00",X"EC",X"D5",X"EC",X"FA",X"EC",X"7F",X"A6",X"70",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"28",X"43",X"29",X"20",X"31",X"39",
		X"38",X"34",X"2C",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",
		X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
