library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity turkey_shoot_bank_a is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of turkey_shoot_bank_a is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"04",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"40",X"04",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"44",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"40",X"04",
		X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"04",X"44",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"44",X"00",X"44",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"04",X"44",X"00",X"00",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"44",X"00",X"44",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"00",X"40",X"04",X"44",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"40",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"40",
		X"04",X"44",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"40",X"04",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"04",X"40",X"04",X"44",X"00",X"04",
		X"40",X"00",X"00",X"00",X"40",X"04",X"40",X"00",X"44",X"40",X"04",X"44",X"00",X"00",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"44",X"00",X"04",X"40",X"04",X"44",X"00",X"04",X"40",X"00",X"00",X"04",
		X"00",X"44",X"40",X"00",X"44",X"00",X"04",X"40",X"00",X"04",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"44",X"40",
		X"44",X"40",X"04",X"00",X"04",X"40",X"00",X"40",X"40",X"00",X"00",X"40",X"00",X"44",X"00",X"04",
		X"44",X"00",X"44",X"40",X"00",X"04",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"40",X"44",X"44",X"44",X"00",
		X"04",X"40",X"00",X"40",X"40",X"00",X"04",X"00",X"00",X"00",X"00",X"04",X"44",X"00",X"44",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"40",X"04",X"44",X"40",X"00",X"04",X"40",X"04",X"00",
		X"40",X"00",X"04",X"00",X"00",X"00",X"00",X"04",X"40",X"00",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"04",X"04",X"40",X"04",X"44",X"00",X"00",X"04",X"40",X"04",X"00",X"40",X"00",X"40",X"00",
		X"00",X"00",X"00",X"44",X"40",X"04",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"04",X"04",X"00",
		X"00",X"00",X"00",X"00",X"04",X"00",X"40",X"04",X"40",X"00",X"40",X"00",X"44",X"40",X"00",X"44",
		X"40",X"04",X"44",X"00",X"04",X"44",X"00",X"00",X"44",X"40",X"44",X"00",X"00",X"44",X"00",X"04",
		X"40",X"00",X"44",X"00",X"00",X"44",X"00",X"00",X"00",X"04",X"00",X"40",X"00",X"00",X"00",X"00",
		X"04",X"00",X"40",X"04",X"40",X"04",X"00",X"04",X"04",X"40",X"04",X"44",X"00",X"04",X"40",X"00",
		X"04",X"44",X"00",X"04",X"40",X"04",X"44",X"00",X"04",X"04",X"40",X"40",X"44",X"04",X"04",X"40",
		X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"00",X"04",
		X"40",X"04",X"00",X"40",X"44",X"00",X"04",X"44",X"00",X"44",X"40",X"00",X"44",X"40",X"00",X"44",
		X"00",X"04",X"40",X"00",X"40",X"04",X"44",X"00",X"44",X"40",X"04",X"40",X"04",X"04",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"40",X"00",X"04",X"40",X"40",X"00",X"00",
		X"44",X"00",X"44",X"40",X"00",X"44",X"40",X"00",X"44",X"40",X"04",X"44",X"00",X"04",X"40",X"00",
		X"40",X"04",X"40",X"04",X"44",X"00",X"44",X"00",X"40",X"04",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"04",X"40",X"40",X"00",X"04",X"40",X"04",X"04",X"40",
		X"04",X"04",X"40",X"04",X"44",X"00",X"04",X"40",X"00",X"44",X"40",X"04",X"00",X"44",X"40",X"04",
		X"44",X"00",X"44",X"00",X"40",X"04",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",
		X"40",X"00",X"00",X"04",X"44",X"00",X"00",X"04",X"40",X"40",X"04",X"40",X"40",X"04",X"40",X"40",
		X"44",X"00",X"04",X"40",X"00",X"44",X"00",X"04",X"00",X"44",X"00",X"04",X"40",X"00",X"44",X"04",
		X"40",X"04",X"44",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",
		X"44",X"00",X"00",X"44",X"00",X"40",X"44",X"00",X"40",X"44",X"00",X"44",X"40",X"00",X"44",X"40",
		X"00",X"44",X"00",X"40",X"00",X"44",X"00",X"04",X"40",X"00",X"40",X"04",X"40",X"04",X"44",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"44",
		X"04",X"00",X"44",X"04",X"00",X"44",X"04",X"04",X"40",X"04",X"04",X"40",X"04",X"04",X"40",X"40",
		X"04",X"40",X"00",X"44",X"00",X"04",X"40",X"40",X"40",X"04",X"44",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"04",X"40",X"00",X"04",X"40",
		X"00",X"04",X"40",X"00",X"44",X"40",X"00",X"44",X"40",X"00",X"44",X"00",X"04",X"40",X"00",X"44",
		X"00",X"04",X"44",X"00",X"04",X"44",X"40",X"00",X"00",X"00",X"00",X"00",X"0A",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",
		X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",
		X"00",X"00",X"00",X"07",X"77",X"77",X"77",X"77",X"70",X"00",X"00",X"00",X"07",X"77",X"77",X"77",
		X"77",X"77",X"70",X"00",X"07",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"77",X"77",X"77",X"77",X"77",X"70",X"00",X"AC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CA",X"A0",X"00",X"00",
		X"0A",X"AC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"AA",X"00",X"00",
		X"00",X"79",X"99",X"99",X"99",X"99",X"97",X"00",X"00",X"00",X"79",X"99",X"99",X"99",X"99",X"99",
		X"70",X"00",X"79",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"97",
		X"77",X"79",X"99",X"99",X"99",X"99",X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"99",X"99",X"99",X"99",X"99",X"97",X"00",X"AC",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AC",X"A0",X"00",X"00",X"0A",X"CA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"CA",X"00",X"00",X"00",X"79",
		X"77",X"77",X"77",X"77",X"97",X"00",X"00",X"07",X"97",X"77",X"77",X"77",X"77",X"79",X"70",X"00",
		X"79",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"99",X"99",X"97",
		X"77",X"77",X"77",X"77",X"97",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"79",X"77",
		X"77",X"77",X"77",X"77",X"97",X"00",X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"79",X"70",X"00",
		X"00",X"07",X"97",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"79",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"90",X"00",X"00",
		X"00",X"00",X"79",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"97",X"00",X"00",X"00",
		X"00",X"07",X"97",X"00",X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"07",
		X"97",X"00",X"07",X"97",X"00",X"00",X"00",X"00",X"07",X"97",X"00",X"00",X"79",X"70",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"97",X"77",X"97",X"00",X"00",X"00",X"00",
		X"07",X"97",X"70",X"00",X"00",X"00",X"00",X"00",X"07",X"79",X"70",X"00",X"00",X"00",X"00",X"79",
		X"70",X"00",X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"07",X"97",X"00",
		X"79",X"70",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"77",X"77",X"79",X"70",X"00",X"00",X"00",X"00",X"79",
		X"77",X"00",X"00",X"00",X"00",X"00",X"77",X"97",X"00",X"00",X"00",X"00",X"07",X"97",X"00",X"00",
		X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"07",X"97",X"07",X"97",X"00",
		X"00",X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"07",X"97",X"00",X"00",X"00",X"00",X"07",X"97",X"70",
		X"00",X"00",X"00",X"07",X"79",X"70",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"AC",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"CA",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"07",X"97",X"79",X"70",X"00",X"00",X"00",
		X"00",X"79",X"70",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"79",X"70",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"79",X"77",X"00",X"00",
		X"00",X"77",X"97",X"00",X"00",X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AC",X"A0",
		X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",
		X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"07",X"97",X"97",X"00",X"00",X"00",X"00",X"07",X"97",
		X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"79",X"70",X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"00",X"07",X"97",X"70",X"00",X"07",X"79",
		X"70",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",
		X"0A",X"CA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",
		X"00",X"79",X"70",X"00",X"00",X"07",X"99",X"70",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",
		X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"07",X"77",X"77",X"77",X"77",X"77",X"77",X"79",X"70",
		X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"79",X"77",X"00",X"77",X"97",X"00",X"00",
		X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"00",X"AC",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"00",
		X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",
		X"00",X"00",X"00",X"0A",X"AA",X"AA",X"A0",X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"79",
		X"70",X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"00",X"00",
		X"79",X"70",X"00",X"00",X"00",X"79",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"70",X"00",X"00",
		X"00",X"07",X"97",X"00",X"00",X"00",X"00",X"07",X"97",X"77",X"79",X"70",X"00",X"00",X"00",X"00",
		X"79",X"70",X"00",X"00",X"00",X"00",X"AA",X"CC",X"CC",X"CC",X"CC",X"CA",X"00",X"00",X"00",X"0A",
		X"CC",X"CC",X"CC",X"CC",X"CA",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",
		X"00",X"AC",X"CC",X"CC",X"CA",X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"79",X"70",X"00",
		X"00",X"07",X"70",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"79",X"70",
		X"00",X"00",X"07",X"97",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"00",X"00",X"00",X"00",X"00",
		X"79",X"70",X"00",X"00",X"00",X"00",X"79",X"77",X"97",X"00",X"00",X"00",X"00",X"07",X"97",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"AA",X"AC",X"A0",X"00",X"00",X"AC",X"AA",X"AA",
		X"AA",X"AA",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"0A",X"CA",
		X"AA",X"AA",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"07",
		X"00",X"00",X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",
		X"07",X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"97",
		X"00",X"00",X"00",X"00",X"07",X"99",X"70",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",
		X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"0A",X"CA",X"00",X"00",
		X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"07",X"97",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"70",X"00",
		X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"AC",X"A0",
		X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"0A",X"CA",X"00",X"00",X"AC",X"A0",
		X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"07",
		X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"07",X"97",X"77",X"77",
		X"77",X"77",X"77",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"97",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",
		X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"0A",X"CA",X"00",X"00",X"AC",X"A0",X"00",X"00",
		X"0A",X"CA",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"70",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"79",X"99",X"99",X"99",X"99",
		X"99",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",
		X"00",X"00",X"0A",X"CA",X"00",X"00",X"0A",X"CA",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",
		X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"07",X"77",X"77",X"77",X"77",X"79",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AC",
		X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",
		X"0A",X"CA",X"00",X"00",X"0A",X"CA",X"AA",X"AA",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",
		X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"07",X"97",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",
		X"00",X"AC",X"A0",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",
		X"00",X"00",X"00",X"AC",X"CC",X"CC",X"CA",X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"79",
		X"70",X"00",X"00",X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",
		X"A0",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",
		X"00",X"0A",X"AA",X"AA",X"A0",X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"79",X"70",X"00",
		X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",
		X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",
		X"00",X"07",X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",
		X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",
		X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"97",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"AC",X"A0",
		X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"07",X"97",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"97",
		X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",
		X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"CA",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"70",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"07",X"77",X"77",X"77",X"77",
		X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"97",X"00",X"00",
		X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",
		X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"CA",
		X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"97",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"79",X"99",X"99",X"99",X"99",X"99",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"79",
		X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AC",
		X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",
		X"0A",X"CA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"CC",X"CC",X"CA",X"00",X"00",
		X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",
		X"00",X"00",X"79",X"70",X"00",X"00",X"07",X"97",X"77",X"77",X"77",X"77",X"77",X"70",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"79",X"70",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",
		X"00",X"AC",X"A0",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",
		X"00",X"00",X"0A",X"AA",X"00",X"00",X"00",X"00",X"0A",X"CA",X"AA",X"AA",X"00",X"00",X"00",X"79",
		X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"00",X"00",X"00",
		X"79",X"70",X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",
		X"A0",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",
		X"0A",X"CC",X"A0",X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"00",X"79",X"70",X"00",
		X"00",X"07",X"70",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"79",X"70",
		X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",
		X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"AA",X"AA",X"AA",X"AA",X"CA",X"00",X"00",X"0A",X"CA",
		X"CA",X"00",X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"07",
		X"97",X"00",X"00",X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",
		X"07",X"97",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",
		X"AC",X"A0",X"00",X"00",X"0A",X"CC",X"CC",X"CC",X"CC",X"A0",X"00",X"00",X"0A",X"CA",X"AC",X"A0",
		X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"07",X"99",X"70",
		X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"79",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"97",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"AC",X"A0",
		X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"0A",X"CA",X"0A",X"CA",X"00",X"00",
		X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"07",X"97",X"97",X"00",X"00",
		X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"07",X"77",X"77",
		X"77",X"77",X"77",X"77",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"97",
		X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",X"00",X"AC",X"A0",X"00",X"00",X"00",
		X"00",X"AC",X"A0",X"00",X"00",X"79",X"70",X"00",X"00",X"07",X"97",X"79",X"70",X"00",X"00",X"00",
		X"00",X"79",X"70",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"97",X"00",X"00",
		X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",X"00",X"0A",X"CA",X"00",X"00",X"00",X"00",X"0A",
		X"CA",X"00",X"00",X"79",X"70",X"00",X"00",X"07",X"97",X"07",X"97",X"00",X"00",X"00",X"00",X"07",
		X"97",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"79",
		X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AC",
		X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"00",X"AC",X"A0",
		X"00",X"79",X"70",X"00",X"00",X"07",X"97",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"79",X"70",
		X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"79",X"70",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",
		X"00",X"AC",X"A0",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"CA",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"00",X"0A",X"CA",X"77",X"79",
		X"70",X"00",X"00",X"07",X"97",X"00",X"07",X"97",X"00",X"00",X"00",X"00",X"07",X"97",X"77",X"77",
		X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",
		X"A0",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"CA",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"00",X"AC",X"77",X"79",X"70",X"00",
		X"00",X"07",X"97",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"79",X"77",X"77",X"79",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",
		X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",
		X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"00",X"0A",X"C9",X"99",X"70",X"00",X"00",X"07",
		X"97",X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"00",X"09",X"99",X"99",X"99",X"70",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"97",X"00",X"00",X"00",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AC",X"AA",X"AA",X"AA",X"AC",X"A0",X"00",X"00",X"00",
		X"AC",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"CA",X"00",X"00",
		X"00",X"00",X"AC",X"AA",X"AA",X"AA",X"AA",X"AA",X"C9",X"99",X"77",X"77",X"77",X"77",X"97",X"00",
		X"00",X"00",X"79",X"77",X"77",X"77",X"77",X"79",X"99",X"99",X"99",X"77",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"97",X"77",X"77",X"77",X"79",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"AC",X"CC",X"CC",X"CC",X"CA",X"A0",X"00",X"00",X"00",X"AC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"AA",X"00",X"00",X"00",X"00",
		X"0A",X"CC",X"CC",X"CC",X"CC",X"CC",X"C7",X"79",X"99",X"99",X"99",X"99",X"97",X"00",X"00",X"00",
		X"07",X"99",X"99",X"99",X"99",X"99",X"77",X"77",X"79",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"99",
		X"99",X"99",X"99",X"99",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"0A",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"77",X"77",X"77",X"77",X"77",X"77",X"70",X"00",X"00",X"00",X"00",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"77",X"77",
		X"77",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"00",X"00",X"00",X"66",X"66",X"66",X"66",X"66",X"00",X"00",X"00",X"00",X"06",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"60",X"00",X"00",X"00",X"00",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"00",X"66",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"E6",X"60",X"00",X"06",X"EE",X"EE",X"EE",X"EE",X"E6",X"60",
		X"00",X"00",X"00",X"66",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"66",X"00",X"00",X"00",X"06",X"6E",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"E6",X"60",X"6E",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"6E",X"60",X"00",X"06",X"E6",
		X"66",X"66",X"66",X"6E",X"60",X"00",X"00",X"00",X"6E",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"E6",X"00",X"00",X"00",X"06",X"E6",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"6E",X"60",X"6E",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6E",X"EE",X"EE",X"EE",X"EE",X"66",X"00",X"00",X"00",
		X"6E",X"60",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"6E",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"66",X"66",X"66",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6E",X"60",
		X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"66",X"66",X"66",
		X"66",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",
		X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",
		X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"EE",X"EE",X"EE",X"EE",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"6E",X"60",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"E6",X"66",X"66",X"66",X"66",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"06",X"E6",X"00",
		X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"6E",X"66",X"66",X"66",X"66",X"E6",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6E",X"60",X"6E",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",
		X"60",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"06",X"E6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6E",X"60",X"6E",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",
		X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",
		X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",
		X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6E",
		X"60",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"6E",X"60",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",
		X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"06",X"E6",X"00",X"00",
		X"00",X"6E",X"60",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6E",X"60",X"6E",X"60",X"00",X"00",X"06",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",
		X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"06",X"E6",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6E",X"60",X"6E",X"60",
		X"00",X"00",X"66",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"66",X"00",X"00",X"00",X"06",X"E6",
		X"00",X"00",X"00",X"6E",X"60",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",
		X"6E",X"60",X"00",X"00",X"00",X"66",X"66",X"66",X"66",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",
		X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"66",X"66",X"66",X"60",X"00",X"00",X"00",X"6E",X"60",
		X"00",X"00",X"06",X"E6",X"66",X"66",X"66",X"66",X"60",X"00",X"00",X"00",X"06",X"66",X"66",X"66",
		X"66",X"6E",X"60",X"6E",X"60",X"00",X"00",X"6E",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"60",
		X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"06",X"E6",X"00",X"00",X"00",
		X"6E",X"60",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"06",X"6E",X"EE",X"EE",X"E6",X"60",X"00",
		X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"66",X"EE",X"EE",X"EE",X"66",
		X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"06",X"6E",X"EE",X"EE",X"EE",X"EE",X"66",X"00",X"00",
		X"00",X"66",X"EE",X"EE",X"EE",X"EE",X"E6",X"60",X"6E",X"60",X"00",X"00",X"6E",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",
		X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"06",X"E6",
		X"66",X"66",X"6E",X"60",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",
		X"6E",X"66",X"66",X"66",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"66",X"66",X"66",
		X"66",X"66",X"E6",X"00",X"00",X"00",X"6E",X"66",X"66",X"66",X"66",X"66",X"00",X"6E",X"60",X"00",
		X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",
		X"00",X"00",X"6E",X"60",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"6E",
		X"60",X"00",X"00",X"06",X"E6",X"00",X"00",X"6E",X"60",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",
		X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",
		X"00",X"00",X"6E",X"60",X"00",X"00",X"6E",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"60",X"00",
		X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"66",X"66",X"66",X"E6",X"00",X"00",X"00",X"6E",
		X"60",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"06",X"E6",X"00",X"00",X"6E",X"60",X"00",X"00",
		X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"06",X"E6",X"00",
		X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",
		X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"66",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"66",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"66",X"EE",X"EE",X"EE",
		X"66",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"06",X"E6",X"00",
		X"00",X"6E",X"60",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",
		X"60",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",
		X"06",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",
		X"00",X"06",X"66",X"66",X"66",X"60",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"6E",X"60",
		X"00",X"00",X"06",X"E6",X"00",X"00",X"6E",X"60",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",
		X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",
		X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",
		X"00",X"06",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6E",X"60",
		X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"06",X"E6",X"00",X"00",X"6E",X"60",X"00",X"00",X"06",
		X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"06",X"E6",X"00",X"00",
		X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",
		X"60",X"00",X"00",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"06",X"E6",X"00",X"00",
		X"6E",X"60",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",
		X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",
		X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"6E",X"60",X"00",
		X"00",X"06",X"E6",X"00",X"00",X"6E",X"60",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",
		X"00",X"00",X"00",X"6E",X"60",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",
		X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",
		X"06",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6E",X"60",X"00",
		X"00",X"00",X"6E",X"60",X"00",X"00",X"06",X"E6",X"00",X"00",X"6E",X"60",X"00",X"00",X"06",X"E6",
		X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"06",X"E6",X"00",X"00",X"00",
		X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",
		X"00",X"00",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"06",X"E6",X"00",X"00",X"6E",
		X"60",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",
		X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",
		X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"6E",X"66",X"66",X"66",X"66",X"66",
		X"66",X"60",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",
		X"66",X"66",X"66",X"60",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",
		X"06",X"E6",X"00",X"00",X"6E",X"60",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",
		X"00",X"00",X"6E",X"60",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"66",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",
		X"E6",X"00",X"00",X"00",X"66",X"EE",X"EE",X"EE",X"66",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",
		X"00",X"6E",X"60",X"00",X"00",X"06",X"E6",X"00",X"00",X"6E",X"60",X"00",X"00",X"06",X"E6",X"00",
		X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",
		X"00",X"00",X"00",X"00",X"06",X"66",X"66",X"66",X"66",X"66",X"66",X"6E",X"60",X"00",X"00",X"06",
		X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"66",X"66",X"66",X"E6",X"00",X"00",
		X"00",X"6E",X"60",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"06",X"E6",X"00",X"00",X"6E",X"60",
		X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"06",
		X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",
		X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"60",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",
		X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"06",
		X"E6",X"00",X"00",X"6E",X"60",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",
		X"00",X"6E",X"60",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"60",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",
		X"00",X"00",X"00",X"6E",X"60",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",
		X"6E",X"60",X"00",X"00",X"06",X"E6",X"00",X"00",X"6E",X"60",X"00",X"00",X"06",X"E6",X"00",X"00",
		X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",
		X"00",X"00",X"00",X"06",X"66",X"66",X"66",X"66",X"66",X"66",X"6E",X"60",X"00",X"00",X"06",X"E6",
		X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"06",X"E6",X"00",X"00",X"00",
		X"6E",X"60",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"06",X"E6",X"66",X"66",X"6E",X"60",X"00",
		X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"66",X"66",X"66",X"E6",
		X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",
		X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"6E",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"E6",
		X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",
		X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"06",X"6E",
		X"EE",X"EE",X"E6",X"60",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",
		X"66",X"EE",X"EE",X"EE",X"66",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"6E",X"66",X"66",
		X"66",X"66",X"66",X"66",X"60",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",
		X"00",X"00",X"6E",X"60",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"6E",
		X"60",X"00",X"00",X"00",X"66",X"66",X"66",X"66",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",
		X"06",X"E6",X"00",X"00",X"00",X"06",X"66",X"66",X"66",X"60",X"00",X"00",X"00",X"6E",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",
		X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",
		X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",
		X"60",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",
		X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"06",
		X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",
		X"00",X"6E",X"60",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"6E",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",
		X"E6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",
		X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",
		X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",
		X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",
		X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",
		X"60",X"00",X"00",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"06",X"E6",
		X"00",X"00",X"00",X"6E",X"60",X"06",X"66",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"66",X"60",X"06",X"E6",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",
		X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",
		X"6E",X"60",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"6E",X"EE",X"60",X"6E",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"06",X"EE",X"E6",X"06",X"E6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",
		X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",
		X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"66",X"EE",
		X"EE",X"E6",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",
		X"6E",X"EE",X"EE",X"66",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",X"00",X"00",X"00",X"6E",X"60",
		X"00",X"00",X"00",X"00",X"00",X"6E",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"E6",X"00",X"00",X"00",X"06",X"E6",X"66",X"66",X"66",X"6E",X"60",X"00",X"06",X"E6",X"66",
		X"66",X"66",X"6E",X"6E",X"66",X"66",X"6E",X"6E",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"E6",X"E6",X"66",X"66",X"E6",X"E6",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"E6",
		X"66",X"66",X"66",X"6E",X"60",X"00",X"00",X"00",X"00",X"00",X"6E",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"66",X"00",X"00",X"00",X"06",X"6E",X"EE",X"EE",X"EE",X"E6",
		X"60",X"00",X"06",X"EE",X"EE",X"EE",X"EE",X"EE",X"E6",X"00",X"00",X"06",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"60",X"00",X"00",X"6E",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"E6",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"6E",X"EE",X"EE",X"EE",X"E6",X"60",X"00",X"00",X"00",X"00",X"00",X"06",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"60",X"00",X"00",X"00",X"00",
		X"66",X"66",X"66",X"66",X"66",X"00",X"00",X"00",X"66",X"66",X"66",X"66",X"66",X"60",X"00",X"00",
		X"00",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"00",
		X"00",X"00",X"06",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"66",X"66",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"28",X"43",X"29",X"20",X"31",X"39",
		X"38",X"34",X"2C",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",
		X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"FF",X"FF",X"FF",
		X"0A",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"AA",X"CC",X"CC",X"CC",X"CA",X"A0",X"00",
		X"00",X"0A",X"AC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"AA",X"00",
		X"00",X"00",X"00",X"0A",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"AA",X"00",
		X"00",X"00",X"00",X"AA",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"AA",X"00",X"AC",X"AA",X"AA",X"AA",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"CA",X"00",X"00",X"00",X"00",X"AC",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"CA",X"A0",X"00",X"00",X"00",X"AC",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"CA",X"00",X"AC",X"A0",X"00",X"00",X"AC",
		X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",
		X"CA",X"00",X"00",X"00",X"0A",X"CA",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",
		X"AC",X"AA",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"CA",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",X"AA",X"AA",X"AA",X"AC",X"AA",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"CA",X"AA",X"AA",X"AA",X"AC",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",X"00",X"AC",X"A0",X"00",
		X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"CA",X"AA",X"AA",X"AA",X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"CA",X"AA",X"AA",X"AA",X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"CA",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",X"00",X"AC",
		X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"CA",X"AA",X"AA",X"AA",X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"CA",X"AA",X"AA",X"AA",X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",
		X"0A",X"CA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",X"AA",X"AA",
		X"AA",X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",X"AA",
		X"AA",X"AA",X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",
		X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"AA",X"AA",
		X"AA",X"AA",X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"AA",
		X"AA",X"AA",X"AA",X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",
		X"00",X"00",X"0A",X"CA",X"00",X"00",X"0A",X"AC",X"CC",X"CC",X"CA",X"A0",X"00",X"00",X"0A",X"CA",
		X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"AC",X"CC",X"CC",X"CA",X"A0",X"00",X"00",X"0A",
		X"CA",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"AC",X"CC",X"CC",X"CC",X"AA",X"00",X"00",
		X"0A",X"CA",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"0A",
		X"CA",X"AA",X"AA",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",
		X"0A",X"CA",X"AA",X"AA",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"AC",X"A0",X"00",
		X"00",X"0A",X"CA",X"AA",X"AA",X"AA",X"CA",X"00",X"00",X"0A",X"CA",X"00",X"AC",X"A0",X"00",X"00",
		X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"0A",X"CA",X"00",X"00",X"AC",X"A0",X"00",X"00",
		X"0A",X"CA",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"AC",X"A0",X"00",
		X"00",X"0A",X"CA",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"0A",X"CA",
		X"00",X"00",X"0A",X"CA",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",
		X"00",X"0A",X"CA",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"AC",X"A0",
		X"00",X"00",X"0A",X"CA",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"AC",
		X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"0A",X"CA",X"00",X"00",X"0A",X"CA",X"00",X"AC",X"A0",
		X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"0A",X"CA",X"00",X"00",X"AC",X"A0",
		X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"AC",
		X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",
		X"0A",X"CA",X"00",X"00",X"0A",X"CA",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",
		X"CA",X"00",X"00",X"0A",X"CA",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",
		X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",
		X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"0A",X"CA",X"00",X"00",X"0A",X"CA",X"00",
		X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"0A",X"CA",X"AA",X"AA",
		X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"AA",
		X"AA",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",
		X"AA",X"AA",X"AA",X"CA",X"00",X"00",X"0A",X"CA",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",
		X"00",X"0A",X"CA",X"00",X"00",X"0A",X"AC",X"CC",X"CC",X"CA",X"A0",X"00",X"00",X"0A",X"CA",X"00",
		X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"AC",X"CC",X"CC",X"CA",X"A0",X"00",X"00",X"0A",X"CA",
		X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"AC",X"CC",X"CC",X"CC",X"AA",X"00",X"00",X"0A",
		X"CA",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"AA",X"AA",X"AA",X"AA",X"CA",X"00",X"00",X"00",X"AA",
		X"AA",X"AA",X"AA",X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",
		X"00",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"AC",X"A0",X"00",X"00",X"AC",
		X"AA",X"AA",X"AA",X"AA",X"CA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",
		X"CA",X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",
		X"CA",X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"CA",X"00",X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"0A",X"CA",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"AC",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",X"00",X"AC",X"A0",X"00",
		X"00",X"AC",X"AA",X"AA",X"AA",X"AA",X"CA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"CA",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"CA",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"AA",X"AA",X"AA",X"AA",X"CA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"AC",
		X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",
		X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",X"00",X"AC",
		X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"AA",X"AA",X"AA",
		X"AA",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",
		X"0A",X"CA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",
		X"00",X"AC",X"A0",X"00",X"00",X"AA",X"CC",X"CC",X"CC",X"CC",X"AA",X"00",X"00",X"0A",X"CA",X"00",
		X"00",X"00",X"AC",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"0A",X"CA",
		X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"AC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"AA",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"AA",
		X"AA",X"AA",X"AA",X"CA",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"AA",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CA",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",
		X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"CA",X"00",X"00",X"0A",X"CA",
		X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"0A",
		X"CA",X"00",X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AC",X"A0",X"00",X"00",
		X"0A",X"CA",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",
		X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"AC",X"A0",X"00",X"00",
		X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",
		X"0A",X"CA",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",
		X"00",X"0A",X"CA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AC",X"A0",
		X"00",X"00",X"0A",X"CA",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"AC",X"A0",
		X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"AC",X"A0",
		X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",
		X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"AA",X"AA",X"AA",X"AA",
		X"CA",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",
		X"AC",X"A0",X"00",X"00",X"AA",X"CC",X"CC",X"CC",X"CC",X"AA",X"00",X"00",X"0A",X"CA",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",
		X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"CA",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"AA",X"AA",
		X"AA",X"AA",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",X"0A",X"CA",X"00",
		X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",
		X"CA",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"CA",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"AC",X"A0",X"00",X"00",X"AC",
		X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",X"0A",
		X"CA",X"00",X"00",X"00",X"AC",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"CA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",
		X"00",X"0A",X"CA",X"00",X"AC",X"A0",X"00",X"00",X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"CA",X"00",X"00",X"0A",X"CA",X"00",X"00",X"00",X"AA",X"CA",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"AC",X"AA",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AC",X"A0",X"00",X"00",X"0A",X"CA",X"00",X"AC",X"AA",X"AA",
		X"AA",X"AC",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"CA",X"AA",
		X"AA",X"AA",X"CA",X"00",X"00",X"00",X"0A",X"AC",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"CA",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AC",
		X"AA",X"AA",X"AA",X"AA",X"CA",X"00",X"AC",X"CC",X"CC",X"CC",X"CA",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"AC",X"CC",X"CC",X"CC",X"AA",X"00",X"00",X"00",X"00",
		X"AA",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CA",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"CC",X"CC",X"CC",X"CC",X"AA",X"00",X"0A",
		X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"F0",X"00",X"0F",X"0F",X"00",X"F0",X"00",X"F0",X"F0",X"00",X"F0",X"FF",X"FF",X"F0",X"F0",
		X"00",X"F0",X"F0",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"0F",X"00",
		X"F0",X"0F",X"00",X"F0",X"0F",X"FF",X"00",X"0F",X"00",X"F0",X"0F",X"00",X"F0",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"0F",X"00",X"F0",X"F0",X"00",X"00",X"F0",
		X"00",X"00",X"F0",X"00",X"00",X"0F",X"00",X"F0",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"00",X"0F",X"00",X"F0",X"0F",X"00",X"F0",X"0F",X"00",X"F0",X"0F",X"00",X"F0",
		X"0F",X"00",X"F0",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"F0",X"0F",
		X"00",X"F0",X"0F",X"0F",X"00",X"0F",X"FF",X"00",X"0F",X"0F",X"00",X"0F",X"00",X"F0",X"FF",X"FF",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"F0",X"0F",X"00",X"F0",X"0F",X"0F",X"00",
		X"0F",X"FF",X"00",X"0F",X"0F",X"00",X"0F",X"00",X"00",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"0F",X"00",X"0F",X"FF",
		X"00",X"F0",X"0F",X"00",X"0F",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"0F",X"00",X"00",X"0F",X"FF",X"00",X"0F",X"00",X"F0",X"0F",X"00",X"F0",X"0F",X"00",X"F0",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",
		X"00",X"F0",X"0F",X"00",X"F0",X"00",X"00",X"F0",X"0F",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",X"0F",X"00",X"0F",X"FF",X"00",X"F0",X"0F",X"00",X"F0",
		X"0F",X"00",X"F0",X"0F",X"00",X"0F",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"FF",X"00",X"F0",X"00",X"F0",X"FF",X"FF",X"00",X"F0",X"00",X"00",
		X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"F0",X"F0",X"00",
		X"F0",X"00",X"0F",X"FF",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",X"0F",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"FF",X"00",X"F0",X"00",X"F0",X"F0",X"00",X"00",X"F0",X"FF",X"F0",
		X"F0",X"00",X"F0",X"F0",X"0F",X"F0",X"0F",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"00",X"F0",X"F0",X"00",X"F0",X"F0",X"00",X"F0",X"FF",X"FF",X"F0",X"F0",X"00",X"F0",X"F0",X"00",
		X"F0",X"F0",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"00",X"00",X"F0",X"00",
		X"00",X"F0",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",X"0F",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",X"0F",X"00",X"00",X"0F",X"00",X"00",X"0F",
		X"00",X"F0",X"0F",X"00",X"F0",X"0F",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"F0",X"F0",X"0F",X"00",X"F0",X"0F",X"0F",X"00",X"0F",X"F0",X"00",X"0F",X"0F",X"00",X"0F",
		X"00",X"F0",X"FF",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",X"0F",X"00",
		X"00",X"0F",X"00",X"00",X"0F",X"00",X"00",X"0F",X"00",X"00",X"0F",X"00",X"F0",X"FF",X"FF",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",X"F0",
		X"0F",X"00",X"0F",X"F0",X"00",X"F0",X"00",X"00",X"FF",X"FF",X"00",X"F0",X"00",X"F0",X"0F",X"FF",
		X"00",X"FF",X"00",X"00",X"0F",X"00",X"00",X"0F",X"F0",X"00",X"0F",X"0F",X"00",X"0F",X"0F",X"00",
		X"0F",X"0F",X"00",X"FF",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"0F",X"F0",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",X"0F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"0F",X"00",X"00",X"0F",X"00",X"00",X"0F",X"00",X"F0",X"0F",X"00",X"F0",X"0F",X"00",X"0F",
		X"F0",X"00",X"FF",X"00",X"00",X"0F",X"00",X"00",X"0F",X"0F",X"00",X"0F",X"F0",X"00",X"0F",X"F0",
		X"00",X"0F",X"0F",X"00",X"FF",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",
		X"00",X"F0",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",X"0F",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",X"0F",X"00",X"00",X"0F",X"00",
		X"00",X"0F",X"00",X"00",X"0F",X"00",X"00",X"0F",X"00",X"F0",X"FF",X"FF",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"00",X"F0",X"0F",X"0F",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"F0",X"F0",X"00",X"F0",X"F0",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"F0",X"0F",X"F0",X"F0",X"0F",X"0F",X"F0",X"0F",X"00",X"F0",X"0F",X"00",X"F0",X"0F",X"00",X"F0",
		X"FF",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"00",X"F0",X"00",X"F0",X"F0",
		X"00",X"F0",X"F0",X"00",X"F0",X"F0",X"00",X"F0",X"F0",X"00",X"F0",X"0F",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"0F",X"00",X"F0",X"0F",X"00",X"F0",X"0F",X"FF",X"00",
		X"0F",X"00",X"00",X"0F",X"00",X"00",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"FF",X"00",X"F0",X"00",X"F0",X"F0",X"00",X"F0",X"F0",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",
		X"F0",X"0F",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"F0",X"00",
		X"00",X"F0",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",X"0F",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"0F",X"00",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",X"0F",X"0F",X"00",X"0F",X"0F",X"00",X"0F",
		X"0F",X"00",X"FF",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"FF",X"00",X"F0",X"00",X"F0",X"F0",X"00",X"F0",X"F0",X"00",X"F0",X"0F",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"0F",
		X"00",X"F0",X"0F",X"00",X"F0",X"0F",X"00",X"F0",X"0F",X"FF",X"00",X"0F",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"F0",X"F0",X"0F",X"00",X"F0",X"0F",X"00",
		X"F0",X"0F",X"00",X"0F",X"FF",X"00",X"00",X"0F",X"00",X"00",X"0F",X"F0",X"FF",X"FF",X"00",X"0F",
		X"00",X"F0",X"0F",X"00",X"F0",X"0F",X"FF",X"00",X"0F",X"0F",X"00",X"0F",X"00",X"F0",X"FF",X"F0",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"00",X"F0",X"00",X"F0",X"F0",X"00",X"00",
		X"0F",X"FF",X"00",X"00",X"00",X"F0",X"F0",X"00",X"F0",X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"00",X"F0",X"00",X"00",X"F0",X"00",X"00",X"F0",
		X"00",X"00",X"F0",X"00",X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"F0",
		X"F0",X"00",X"F0",X"F0",X"00",X"F0",X"F0",X"00",X"F0",X"F0",X"00",X"F0",X"F0",X"00",X"F0",X"0F",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"F0",X"F0",X"00",X"F0",X"F0",X"00",
		X"F0",X"F0",X"00",X"F0",X"0F",X"0F",X"00",X"0F",X"0F",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"00",X"F0",X"F0",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"0F",X"0F",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"FF",X"00",X"0F",X"00",X"F0",X"0F",X"00",X"00",X"0F",X"00",X"00",
		X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"0F",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"0F",X"00",X"00",X"FF",X"F0",X"00",X"0F",X"00",X"00",
		X"0F",X"00",X"00",X"0F",X"0F",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"0F",X"F0",X"0F",X"0F",X"00",X"0F",X"0F",X"00",X"0F",X"0F",
		X"00",X"0F",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"0F",X"F0",X"0F",X"0F",X"00",X"0F",X"0F",X"00",X"0F",X"0F",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"F0",X"F0",X"00",X"F0",X"0F",X"0F",X"00",X"00",X"F0",X"00",X"0F",X"0F",X"00",X"F0",
		X"00",X"F0",X"F0",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"F0",X"0F",X"0F",
		X"00",X"0F",X"0F",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",X"0F",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"F0",X"F0",X"00",X"F0",X"00",X"0F",X"00",X"00",
		X"F0",X"00",X"0F",X"00",X"00",X"F0",X"00",X"F0",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"F0",X"0F",X"0F",X"00",X"00",X"F0",X"00",
		X"0F",X"0F",X"00",X"F0",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"0F",X"F0",X"0F",X"0F",X"00",X"0F",X"0F",X"00",X"0F",X"0F",X"00",X"00",X"FF",
		X"00",X"F0",X"0F",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"F0",
		X"F0",X"0F",X"00",X"00",X"F0",X"00",X"0F",X"00",X"F0",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"F0",X"00",X"0F",X"F0",X"00",X"0F",X"F0",X"00",X"0F",X"F0",X"00",X"0F",X"F0",
		X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",
		X"0F",X"0F",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",X"FF",X"FF",
		X"F0",X"0F",X"0F",X"00",X"FF",X"FF",X"F0",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"00",X"0F",X"FF",X"00",X"F0",X"00",X"00",X"0F",X"FF",X"00",X"00",
		X"00",X"F0",X"0F",X"FF",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"F0",X"FF",X"00",X"F0",X"00",X"0F",X"00",X"00",X"F0",X"00",X"0F",X"00",X"00",X"F0",X"0F",X"F0",
		X"F0",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",X"0F",X"0F",X"00",X"00",
		X"F0",X"00",X"0F",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"0F",X"00",X"0F",X"F0",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"0F",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"0F",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",X"0F",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",X"F0",X"F0",
		X"F0",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",X"FF",X"FF",X"F0",X"00",X"F0",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"0F",X"00",
		X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"F0",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"00",X"0F",X"00",X"00",X"F0",X"00",X"0F",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"00",X"F0",X"00",X"F0",X"F0",X"00",X"F0",
		X"F0",X"00",X"F0",X"F0",X"00",X"F0",X"F0",X"00",X"F0",X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"00",X"0F",X"F0",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",X"00",X"F0",
		X"00",X"00",X"F0",X"00",X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",
		X"F0",X"0F",X"00",X"00",X"0F",X"00",X"00",X"F0",X"00",X"0F",X"00",X"00",X"F0",X"00",X"00",X"FF",
		X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"F0",X"F0",X"00",X"F0",X"00",X"0F",
		X"00",X"00",X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"00",X"F0",X"0F",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"FF",X"00",X"0F",X"0F",X"00",X"FF",X"FF",X"F0",X"00",
		X"0F",X"00",X"00",X"0F",X"00",X"00",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"F0",X"00",X"00",X"FF",X"FF",X"00",X"F0",X"00",X"F0",X"00",X"00",X"F0",X"F0",X"00",X"F0",
		X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"00",X"F0",X"00",X"00",X"F0",
		X"FF",X"00",X"FF",X"00",X"F0",X"F0",X"00",X"F0",X"F0",X"00",X"F0",X"0F",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"F0",X"F0",X"00",X"F0",X"00",X"00",X"F0",X"00",X"0F",X"00",
		X"00",X"0F",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"FF",X"00",X"F0",X"00",X"F0",X"F0",X"00",X"F0",X"0F",X"FF",X"00",X"F0",X"00",X"F0",X"F0",X"00",
		X"F0",X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"00",X"F0",X"00",X"F0",
		X"F0",X"00",X"F0",X"0F",X"FF",X"F0",X"00",X"00",X"F0",X"F0",X"00",X"F0",X"0F",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",X"0F",X"F0",X"00",X"00",X"00",
		X"00",X"0F",X"F0",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"F0",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",
		X"F0",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"F0",
		X"00",X"0F",X"00",X"00",X"F0",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"00",X"00",
		X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"0F",X"00",
		X"00",X"F0",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"00",X"F0",
		X"00",X"F0",X"00",X"00",X"F0",X"00",X"FF",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"0F",X"00",X"F0",X"F0",X"0F",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"FF",X"F0",X"F0",X"00",X"00",X"0F",X"FF",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",
		X"F0",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",X"00",X"FF",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",
		X"00",X"F0",X"00",X"00",X"F0",X"00",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"0F",X"00",X"FF",X"FF",X"F0",X"00",X"0F",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"0F",
		X"00",X"00",X"FF",X"FF",X"F0",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"00",X"F0",X"F0",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"00",
		X"F0",X"F0",X"FF",X"00",X"F0",X"F0",X"FF",X"F0",X"0F",X"F0",X"F0",X"00",X"F0",X"00",X"F0",X"00",
		X"0F",X"F0",X"FF",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"00",X"FF",X"F0",X"F0",X"00",
		X"FF",X"00",X"F0",X"00",X"FF",X"F0",X"FF",X"F0",X"F0",X"00",X"FF",X"00",X"F0",X"00",X"F0",X"00",
		X"0F",X"F0",X"F0",X"00",X"FF",X"F0",X"F0",X"F0",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"FF",X"F0",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"FF",X"F0",X"00",X"F0",
		X"00",X"F0",X"00",X"F0",X"F0",X"F0",X"0F",X"00",X"F0",X"00",X"F0",X"F0",X"FF",X"00",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"FF",X"F0",X"F0",X"F0",X"FF",X"F0",
		X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"F0",X"FF",X"00",X"F0",X"F0",X"FF",X"00",
		X"F0",X"00",X"F0",X"00",X"0F",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"F0",X"FF",X"00",
		X"F0",X"F0",X"FF",X"00",X"F0",X"F0",X"F0",X"F0",X"FF",X"F0",X"F0",X"00",X"FF",X"F0",X"00",X"F0",
		X"FF",X"F0",X"FF",X"F0",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"00",
		X"F0",X"F0",X"F0",X"F0",X"FF",X"F0",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"FF",X"F0",
		X"00",X"F0",X"0F",X"00",X"F0",X"00",X"FF",X"F0",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"00",X"00",
		X"0F",X"00",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"FF",X"F0",
		X"FF",X"F0",X"0F",X"00",X"00",X"00",X"0F",X"00",X"F0",X"00",X"0F",X"00",X"00",X"F0",X"0F",X"00",
		X"F0",X"00",X"00",X"F0",X"0F",X"00",X"F0",X"00",X"00",X"F0",X"F0",X"00",X"FF",X"00",X"0F",X"00",
		X"F0",X"F0",X"FF",X"00",X"F0",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",
		X"F0",X"00",X"F0",X"00",X"F0",X"00",X"0F",X"00",X"0F",X"00",X"00",X"F0",X"00",X"F0",X"00",X"F0",
		X"0F",X"00",X"00",X"00",X"0F",X"00",X"F0",X"F0",X"0F",X"00",X"00",X"00",X"0F",X"00",X"0F",X"00",
		X"FF",X"F0",X"0F",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"0F",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"0F",X"00",X"F0",X"00",X"0F",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"00",X"0F",X"00",X"FF",X"00",X"0F",X"00",X"0F",X"00",
		X"FF",X"F0",X"0F",X"00",X"F0",X"F0",X"00",X"F0",X"0F",X"00",X"FF",X"F0",X"FF",X"F0",X"00",X"F0",
		X"FF",X"F0",X"00",X"F0",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"F0",X"00",X"F0",X"00",X"F0",
		X"FF",X"F0",X"FF",X"00",X"00",X"F0",X"00",X"F0",X"FF",X"F0",X"0F",X"F0",X"F0",X"00",X"FF",X"F0",
		X"F0",X"F0",X"FF",X"F0",X"FF",X"F0",X"00",X"F0",X"0F",X"00",X"F0",X"00",X"F0",X"00",X"FF",X"F0",
		X"F0",X"F0",X"FF",X"F0",X"F0",X"F0",X"FF",X"F0",X"FF",X"F0",X"F0",X"F0",X"FF",X"F0",X"00",X"F0",
		X"00",X"F0",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"0F",X"00",X"F0",X"00",X"00",X"F0",X"0F",X"00",X"F0",X"00",X"0F",X"00",X"00",X"F0",
		X"00",X"00",X"FF",X"F0",X"00",X"00",X"FF",X"F0",X"00",X"00",X"F0",X"00",X"0F",X"00",X"00",X"F0",
		X"0F",X"00",X"F0",X"00",X"0F",X"00",X"F0",X"F0",X"00",X"F0",X"0F",X"00",X"0F",X"00",X"0F",X"00",
		X"FF",X"F0",X"F0",X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",
		X"0F",X"00",X"00",X"F0",X"00",X"00",X"0F",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"0F",X"F0",
		X"00",X"00",X"0F",X"00",X"0F",X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"FF",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",
		X"54",X"20",X"28",X"43",X"29",X"20",X"31",X"39",X"38",X"34",X"2C",X"20",X"57",X"49",X"4C",X"4C",
		X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",
		X"20",X"49",X"4E",X"43",X"2E",X"DD",X"DD",X"D0",X"DD",X"DD",X"D0",X"DD",X"DD",X"D0",X"DD",X"DD",
		X"D0",X"DD",X"DD",X"D0",X"DD",X"DD",X"D0",X"DD",X"DD",X"D0",X"DD",X"DD",X"D0",X"DD",X"DD",X"D0",
		X"DD",X"D0",X"DD",X"D0",X"DD",X"D0",X"DD",X"D0",X"DD",X"D0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
