library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity turkey_shoot_prog2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of turkey_shoot_prog2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"28",X"43",X"29",X"20",X"31",X"39",
		X"38",X"34",X"2C",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",
		X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"34",X"06",X"B7",
		X"CB",X"00",X"97",X"85",X"C6",X"20",X"3D",X"C3",X"80",X"00",X"DD",X"86",X"35",X"86",X"34",X"06",
		X"B7",X"CB",X"20",X"97",X"88",X"C6",X"20",X"3D",X"C3",X"80",X"00",X"DD",X"89",X"35",X"86",X"34",
		X"04",X"F6",X"CB",X"E0",X"C1",X"F8",X"23",X"F9",X"35",X"84",X"34",X"51",X"1A",X"50",X"8D",X"EF",
		X"1F",X"01",X"DE",X"86",X"CC",X"03",X"10",X"B7",X"C8",X"00",X"AF",X"C1",X"5A",X"26",X"FB",X"86",
		X"06",X"B7",X"C8",X"00",X"35",X"D1",X"34",X"51",X"1A",X"50",X"8D",X"D3",X"5F",X"48",X"CE",X"E3",
		X"00",X"EE",X"C6",X"10",X"9E",X"86",X"34",X"40",X"8D",X"0A",X"35",X"40",X"10",X"8E",X"AD",X"ED",
		X"8D",X"0F",X"35",X"D1",X"C6",X"03",X"F7",X"C8",X"00",X"8D",X"06",X"C6",X"06",X"F7",X"C8",X"00",
		X"39",X"34",X"1F",X"1A",X"50",X"1F",X"41",X"32",X"25",X"37",X"2E",X"34",X"2E",X"32",X"6A",X"37",
		X"2E",X"34",X"2E",X"32",X"6A",X"37",X"2E",X"34",X"2E",X"32",X"6A",X"37",X"2E",X"34",X"2E",X"32",
		X"6A",X"37",X"2E",X"34",X"2E",X"32",X"6A",X"37",X"2E",X"34",X"2E",X"32",X"67",X"37",X"20",X"34",
		X"20",X"31",X"62",X"1F",X"14",X"35",X"9F",X"34",X"01",X"1A",X"50",X"CE",X"AD",X"ED",X"10",X"9E",
		X"86",X"8D",X"B1",X"35",X"81",X"BD",X"DF",X"C4",X"4F",X"BD",X"66",X"BC",X"4F",X"8D",X"87",X"4F",
		X"34",X"01",X"1A",X"50",X"BD",X"DF",X"C4",X"B7",X"C8",X"81",X"CC",X"00",X"00",X"FD",X"C8",X"84",
		X"CC",X"C0",X"C0",X"FD",X"C8",X"86",X"86",X"10",X"B7",X"C8",X"80",X"BD",X"DF",X"C4",X"35",X"81",
		X"34",X"07",X"1A",X"50",X"BD",X"E0",X"4F",X"86",X"03",X"B7",X"C8",X"00",X"DC",X"89",X"FD",X"C8",
		X"84",X"CC",X"08",X"20",X"FD",X"C8",X"86",X"7F",X"C8",X"81",X"86",X"10",X"B7",X"C8",X"80",X"BD",
		X"DF",X"C4",X"86",X"06",X"B7",X"C8",X"00",X"35",X"87",X"7A",X"AE",X"5B",X"2E",X"32",X"C6",X"03",
		X"F7",X"C8",X"00",X"86",X"04",X"B7",X"AE",X"5B",X"BE",X"AE",X"59",X"EC",X"84",X"26",X"05",X"8E",
		X"E2",X"DE",X"EC",X"84",X"FD",X"80",X"16",X"EC",X"02",X"FD",X"80",X"18",X"EC",X"04",X"FD",X"80",
		X"1A",X"EC",X"06",X"FD",X"80",X"1C",X"30",X"08",X"BF",X"AE",X"59",X"86",X"06",X"B7",X"C8",X"00",
		X"8D",X"01",X"39",X"7A",X"AE",X"57",X"2E",X"32",X"C6",X"03",X"F7",X"C8",X"00",X"86",X"03",X"B7",
		X"AE",X"57",X"BE",X"AE",X"55",X"EC",X"84",X"26",X"05",X"8E",X"E2",X"C4",X"EC",X"84",X"FD",X"80",
		X"0E",X"EC",X"02",X"FD",X"80",X"10",X"EC",X"04",X"FD",X"80",X"12",X"EC",X"06",X"FD",X"80",X"14",
		X"30",X"08",X"BF",X"AE",X"55",X"86",X"06",X"B7",X"C8",X"00",X"39",X"C6",X"03",X"F7",X"C8",X"00",
		X"7A",X"AE",X"51",X"2E",X"23",X"86",X"04",X"B7",X"AE",X"51",X"BE",X"AE",X"4F",X"EC",X"84",X"26",
		X"05",X"8E",X"E2",X"9C",X"EC",X"84",X"FD",X"87",X"86",X"EC",X"02",X"FD",X"87",X"88",X"EC",X"04",
		X"FD",X"87",X"8A",X"30",X"06",X"BF",X"AE",X"4F",X"7A",X"AE",X"54",X"2E",X"23",X"86",X"09",X"B7",
		X"AE",X"54",X"BE",X"AE",X"52",X"EC",X"84",X"26",X"05",X"8E",X"E2",X"B0",X"EC",X"84",X"FD",X"87",
		X"82",X"EC",X"02",X"FD",X"87",X"80",X"EC",X"04",X"FD",X"87",X"96",X"30",X"06",X"BF",X"AE",X"52",
		X"86",X"06",X"B7",X"C8",X"00",X"39",X"CE",X"E2",X"34",X"96",X"09",X"27",X"03",X"CE",X"E2",X"40",
		X"37",X"36",X"A7",X"84",X"E7",X"A4",X"37",X"36",X"A7",X"84",X"E7",X"A4",X"8E",X"E2",X"B0",X"BF",
		X"AE",X"52",X"8E",X"E2",X"58",X"BF",X"AE",X"4F",X"39",X"CE",X"E2",X"4C",X"7F",X"AE",X"51",X"7F",
		X"AE",X"54",X"20",X"DC",X"A5",X"A4",X"C0",X"B9",X"C0",X"A9",X"50",X"4F",X"C0",X"09",X"C0",X"19",
		X"25",X"24",X"C0",X"09",X"C0",X"19",X"D0",X"CF",X"C0",X"B9",X"C0",X"A9",X"25",X"24",X"C0",X"09",
		X"C0",X"19",X"A5",X"A4",X"C0",X"B9",X"C0",X"A9",X"0F",X"F0",X"F0",X"F0",X"00",X"FF",X"F0",X"D0",
		X"00",X"DF",X"0F",X"D0",X"00",X"CF",X"0F",X"C0",X"F0",X"C0",X"0F",X"B0",X"F0",X"B0",X"00",X"BF",
		X"F0",X"A0",X"00",X"AF",X"0F",X"A0",X"00",X"9F",X"0F",X"90",X"F0",X"90",X"0F",X"80",X"F0",X"80",
		X"00",X"8F",X"F0",X"70",X"00",X"7F",X"0F",X"70",X"00",X"6F",X"0F",X"60",X"F0",X"60",X"0F",X"50",
		X"F0",X"50",X"00",X"5F",X"F0",X"40",X"00",X"4F",X"0F",X"40",X"00",X"00",X"1E",X"80",X"2F",X"00",
		X"2F",X"40",X"2F",X"00",X"2F",X"40",X"1E",X"80",X"2F",X"40",X"1E",X"80",X"2F",X"00",X"00",X"00",
		X"DF",X"D9",X"0F",X"D6",X"0F",X"D6",X"0F",X"D6",X"DF",X"D9",X"0F",X"D6",X"0F",X"D6",X"0F",X"D6",
		X"DF",X"D9",X"00",X"00",X"0D",X"ED",X"0A",X"EE",X"0F",X"EA",X"00",X"00",X"0A",X"EE",X"0F",X"EA",
		X"0D",X"ED",X"00",X"00",X"0F",X"EA",X"0D",X"ED",X"0A",X"EE",X"00",X"00",X"00",X"00",X"FF",X"FA",
		X"FF",X"8A",X"FF",X"BA",X"FF",X"DA",X"FF",X"DA",X"FF",X"FA",X"FF",X"8A",X"FF",X"BA",X"FF",X"BA",
		X"FF",X"DA",X"FF",X"FA",X"FF",X"8A",X"FF",X"8A",X"FF",X"BA",X"FF",X"DA",X"FF",X"FA",X"00",X"00",
		X"E3",X"0E",X"E3",X"2E",X"E3",X"4E",X"E3",X"6E",X"E3",X"8E",X"E3",X"AE",X"E3",X"CE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"EE",X"F0",X"BF",X"FF",X"1F",X"D2",X"1E",X"B0",X"B7",X"ED",X"AE",X"E9",X"01",X"FE",
		X"01",X"DD",X"01",X"BD",X"AF",X"E1",X"97",X"EA",X"FF",X"BE",X"2F",X"50",X"00",X"00",X"00",X"00",
		X"FF",X"EF",X"FF",X"EF",X"BF",X"CF",X"EF",X"EB",X"CF",X"FA",X"AE",X"DF",X"D6",X"FE",X"FF",X"6F",
		X"FF",X"AF",X"4F",X"F1",X"FF",X"6F",X"DF",X"F1",X"FF",X"FF",X"E6",X"FF",X"0F",X"F0",X"00",X"00",
		X"FF",X"F0",X"0F",X"FF",X"FF",X"F0",X"AF",X"E1",X"F0",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"F0",X"0F",X"F0",X"F0",X"D0",X"00",X"00",X"00",X"FF",X"00",X"00",X"0F",X"C0",
		X"F0",X"C0",X"00",X"CF",X"FF",X"CF",X"FF",X"C0",X"F0",X"CF",X"0F",X"CF",X"00",X"00",X"0F",X"C0",
		X"0F",X"C0",X"F0",X"C0",X"F0",X"C0",X"00",X"CF",X"00",X"CF",X"00",X"00",X"00",X"00",X"FF",X"CF",
		X"FF",X"CF",X"FF",X"C0",X"FF",X"C0",X"F0",X"CF",X"F0",X"CF",X"0F",X"CF",X"0F",X"CF",X"00",X"00",
		X"0F",X"FF",X"F0",X"FF",X"FF",X"F0",X"FF",X"FF",X"00",X"FF",X"F0",X"F0",X"0F",X"F0",X"0F",X"FF",
		X"0F",X"F0",X"F0",X"F0",X"00",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"FF",X"0F",X"FF",X"A6",X"C4",
		X"2D",X"2D",X"34",X"40",X"CE",X"AE",X"2D",X"48",X"AE",X"C6",X"30",X"1F",X"AF",X"C6",X"26",X"19",
		X"10",X"8E",X"AE",X"0D",X"AE",X"A6",X"AE",X"04",X"AF",X"A6",X"10",X"AE",X"02",X"10",X"AF",X"C6",
		X"10",X"AE",X"00",X"8E",X"AD",X"ED",X"10",X"AF",X"86",X"35",X"40",X"33",X"43",X"20",X"CF",X"39",
		X"A6",X"C4",X"2D",X"17",X"8E",X"AE",X"0D",X"48",X"10",X"AE",X"41",X"10",X"AF",X"86",X"8E",X"AE",
		X"2D",X"10",X"AE",X"22",X"10",X"AF",X"86",X"33",X"43",X"20",X"E5",X"39",X"BD",X"00",X"3F",X"F6",
		X"C9",X"85",X"2A",X"3D",X"CC",X"35",X"3D",X"F7",X"C9",X"85",X"F6",X"C9",X"84",X"B7",X"C9",X"85",
		X"B6",X"C9",X"84",X"88",X"80",X"0D",X"28",X"26",X"02",X"DD",X"4E",X"AD",X"9F",X"BF",X"33",X"BD",
		X"6F",X"E9",X"86",X"14",X"B7",X"C9",X"00",X"D6",X"47",X"27",X"02",X"0A",X"47",X"D6",X"8D",X"26",
		X"0C",X"03",X"8D",X"B6",X"C9",X"87",X"2B",X"10",X"CC",X"E4",X"8B",X"DD",X"35",X"BD",X"00",X"4E",
		X"3B",X"B6",X"C9",X"86",X"6E",X"9F",X"BF",X"35",X"B6",X"C9",X"86",X"97",X"50",X"0F",X"5D",X"DC",
		X"2F",X"2A",X"20",X"86",X"FF",X"90",X"94",X"97",X"92",X"BD",X"F6",X"A3",X"BD",X"F6",X"B6",X"96",
		X"29",X"2A",X"06",X"BD",X"EC",X"4D",X"BD",X"EC",X"5A",X"DC",X"2D",X"DD",X"2F",X"96",X"28",X"26",
		X"02",X"03",X"28",X"B6",X"CB",X"E0",X"97",X"94",X"BD",X"F6",X"DC",X"BD",X"F6",X"C9",X"B6",X"CB",
		X"E0",X"90",X"94",X"97",X"94",X"B6",X"CB",X"E0",X"81",X"80",X"22",X"0E",X"CC",X"E4",X"D3",X"DD",
		X"35",X"20",X"48",X"CC",X"E4",X"DD",X"DD",X"35",X"20",X"41",X"B6",X"C9",X"86",X"BD",X"F9",X"59",
		X"26",X"03",X"BD",X"F9",X"CD",X"DC",X"2F",X"83",X"00",X"01",X"DD",X"2F",X"2A",X"0F",X"86",X"7F",
		X"90",X"93",X"97",X"91",X"BD",X"00",X"5A",X"BD",X"F6",X"99",X"BD",X"F6",X"AC",X"B6",X"CB",X"E0",
		X"97",X"93",X"BD",X"F6",X"D2",X"BD",X"F6",X"BF",X"B6",X"CB",X"E0",X"90",X"93",X"97",X"93",X"CC",
		X"E5",X"18",X"DD",X"35",X"0F",X"8D",X"20",X"03",X"B6",X"C9",X"86",X"BD",X"00",X"4E",X"3B",X"BD",
		X"27",X"6F",X"0F",X"28",X"BD",X"00",X"48",X"BD",X"3E",X"78",X"0D",X"28",X"27",X"FC",X"BD",X"00",
		X"39",X"39",X"34",X"01",X"1A",X"50",X"C6",X"00",X"BD",X"E5",X"61",X"20",X"04",X"34",X"01",X"1A",
		X"50",X"CC",X"E5",X"18",X"DD",X"35",X"0F",X"8D",X"BD",X"DF",X"81",X"BD",X"FA",X"10",X"BD",X"7E",
		X"56",X"35",X"81",X"DE",X"48",X"AE",X"C3",X"26",X"04",X"DE",X"4A",X"AE",X"C3",X"DF",X"48",X"6E",
		X"84",X"34",X"01",X"1A",X"50",X"D7",X"29",X"8E",X"E5",X"76",X"AE",X"85",X"9F",X"33",X"9F",X"4A",
		X"9F",X"48",X"35",X"81",X"E5",X"A5",X"E5",X"86",X"E5",X"D7",X"E5",X"FF",X"E6",X"2A",X"E6",X"4F",
		X"E6",X"81",X"E6",X"9D",X"E6",X"A7",X"BD",X"E7",X"03",X"BD",X"F5",X"FD",X"BD",X"00",X"DE",X"BD",
		X"E6",X"5F",X"39",X"00",X"00",X"ED",X"A5",X"34",X"56",X"E6",X"5F",X"65",X"A5",X"01",X"0C",X"66",
		X"69",X"66",X"55",X"D5",X"F5",X"B6",X"CB",X"E0",X"81",X"F0",X"25",X"0C",X"BD",X"E7",X"03",X"BD",
		X"D1",X"17",X"BD",X"E1",X"AB",X"BD",X"F5",X"FD",X"BD",X"E5",X"53",X"BD",X"00",X"DE",X"BD",X"7E",
		X"D6",X"BD",X"D5",X"4B",X"39",X"00",X"00",X"E6",X"67",X"E6",X"5F",X"D5",X"F5",X"D5",X"A1",X"E5",
		X"92",X"E5",X"92",X"E5",X"92",X"E5",X"92",X"BD",X"E7",X"03",X"BD",X"E0",X"D7",X"BD",X"F5",X"FD",
		X"BD",X"01",X"29",X"BD",X"00",X"DE",X"BD",X"E5",X"53",X"BD",X"D5",X"4B",X"39",X"00",X"00",X"E6",
		X"5F",X"D5",X"F5",X"D5",X"A7",X"66",X"5D",X"66",X"4D",X"E5",X"92",X"E5",X"92",X"E5",X"92",X"BD",
		X"E7",X"03",X"BD",X"F5",X"FD",X"BD",X"13",X"21",X"BD",X"01",X"29",X"BD",X"00",X"DE",X"BD",X"E5",
		X"53",X"BD",X"DD",X"82",X"BD",X"D5",X"4B",X"39",X"00",X"00",X"E6",X"67",X"E6",X"5F",X"D5",X"F5",
		X"D5",X"AD",X"E5",X"92",X"E5",X"92",X"E5",X"92",X"E5",X"92",X"BD",X"E7",X"03",X"BD",X"E1",X"73",
		X"BD",X"01",X"29",X"BD",X"00",X"DE",X"BD",X"E5",X"53",X"BD",X"D5",X"4B",X"39",X"00",X"00",X"E6",
		X"5F",X"D5",X"F5",X"D5",X"AD",X"E5",X"92",X"E5",X"92",X"E5",X"92",X"E5",X"92",X"E5",X"92",X"BD",
		X"01",X"29",X"BD",X"E1",X"39",X"BD",X"00",X"DE",X"BD",X"E5",X"53",X"BD",X"D5",X"4B",X"39",X"96",
		X"60",X"27",X"03",X"7E",X"F1",X"CA",X"39",X"96",X"47",X"27",X"03",X"7E",X"D5",X"09",X"39",X"00",
		X"00",X"D5",X"B3",X"E5",X"92",X"E5",X"92",X"E5",X"92",X"E5",X"92",X"E5",X"92",X"E5",X"92",X"E5",
		X"92",X"BD",X"D5",X"86",X"BD",X"00",X"DE",X"BD",X"E5",X"53",X"39",X"00",X"00",X"D5",X"B3",X"E5",
		X"92",X"E5",X"92",X"E5",X"92",X"E5",X"92",X"E5",X"92",X"E5",X"92",X"E5",X"92",X"BD",X"D5",X"86",
		X"BD",X"00",X"DE",X"BD",X"E5",X"53",X"39",X"BD",X"D5",X"86",X"39",X"34",X"71",X"1A",X"50",X"CC",
		X"03",X"03",X"9E",X"89",X"FE",X"C5",X"83",X"20",X"07",X"34",X"71",X"1A",X"50",X"CC",X"06",X"05",
		X"BD",X"E0",X"4F",X"7F",X"CB",X"A0",X"F7",X"C8",X"00",X"10",X"8E",X"BC",X"DD",X"F6",X"C5",X"82",
		X"27",X"17",X"C6",X"40",X"BD",X"DF",X"CD",X"BD",X"E0",X"4F",X"10",X"8E",X"BD",X"5D",X"30",X"89",
		X"00",X"80",X"BD",X"DF",X"CD",X"10",X"8E",X"BD",X"DD",X"B7",X"C8",X"00",X"F6",X"C5",X"81",X"27",
		X"07",X"37",X"10",X"AF",X"A1",X"5A",X"26",X"F9",X"CC",X"06",X"01",X"B7",X"C8",X"00",X"F7",X"CB",
		X"A0",X"35",X"F1",X"96",X"A9",X"27",X"27",X"86",X"03",X"B7",X"C8",X"00",X"8E",X"BC",X"DD",X"F6",
		X"C5",X"82",X"27",X"09",X"10",X"9E",X"89",X"BD",X"DF",X"D3",X"8E",X"BD",X"DD",X"F6",X"C5",X"81",
		X"27",X"07",X"10",X"BE",X"C5",X"83",X"BD",X"DF",X"D3",X"86",X"06",X"B7",X"C8",X"00",X"39",X"BD",
		X"E5",X"1F",X"5F",X"BD",X"E5",X"61",X"BD",X"F0",X"6B",X"BD",X"E7",X"FF",X"96",X"25",X"9A",X"26",
		X"27",X"25",X"BD",X"DB",X"1C",X"86",X"FF",X"97",X"9F",X"8D",X"21",X"BD",X"E8",X"5A",X"BD",X"E8",
		X"27",X"BD",X"7E",X"73",X"96",X"25",X"9A",X"26",X"27",X"0A",X"8D",X"10",X"BD",X"E8",X"63",X"BD",
		X"E7",X"FF",X"20",X"03",X"BD",X"7E",X"73",X"86",X"FF",X"97",X"97",X"39",X"BD",X"E9",X"A3",X"BD",
		X"E5",X"1F",X"BD",X"E8",X"CC",X"F1",X"A6",X"7B",X"27",X"20",X"86",X"05",X"BD",X"70",X"08",X"CE",
		X"EC",X"21",X"BD",X"E9",X"37",X"BD",X"E5",X"1F",X"F6",X"A6",X"7A",X"F7",X"A6",X"7B",X"CE",X"EC",
		X"37",X"BD",X"E9",X"37",X"BD",X"E5",X"1F",X"BD",X"E9",X"8D",X"96",X"41",X"85",X"04",X"27",X"4A",
		X"BD",X"00",X"82",X"86",X"01",X"BD",X"70",X"08",X"B6",X"A6",X"7B",X"81",X"1B",X"26",X"02",X"20",
		X"44",X"81",X"17",X"26",X"1C",X"DE",X"23",X"E6",X"5F",X"27",X"2F",X"BD",X"E9",X"62",X"5A",X"E7",
		X"5F",X"A6",X"C5",X"B7",X"A6",X"74",X"CC",X"FF",X"F5",X"BD",X"E9",X"71",X"BD",X"E9",X"8D",X"20",
		X"19",X"DE",X"23",X"E6",X"5F",X"B6",X"A6",X"74",X"A7",X"C5",X"5C",X"E7",X"5F",X"E1",X"5E",X"24",
		X"CE",X"CC",X"00",X"0B",X"BD",X"E9",X"71",X"BD",X"E9",X"66",X"DC",X"55",X"C3",X"FF",X"FF",X"DD",
		X"55",X"10",X"2E",X"FF",X"7A",X"BD",X"E5",X"1F",X"96",X"63",X"9A",X"64",X"26",X"F7",X"39",X"C6",
		X"01",X"CE",X"BB",X"BC",X"8D",X"3E",X"26",X"03",X"BD",X"7E",X"73",X"CE",X"AA",X"27",X"C6",X"0A",
		X"8D",X"32",X"27",X"13",X"D7",X"25",X"C1",X"01",X"27",X"0D",X"BD",X"7E",X"73",X"8D",X"25",X"5A",
		X"2F",X"02",X"D7",X"25",X"BD",X"7E",X"73",X"CE",X"A9",X"48",X"C6",X"25",X"8D",X"16",X"27",X"13",
		X"D7",X"26",X"C1",X"01",X"27",X"0D",X"BD",X"7E",X"73",X"8D",X"09",X"5A",X"2F",X"02",X"D7",X"26",
		X"BD",X"7E",X"73",X"39",X"9E",X"03",X"96",X"05",X"AC",X"C4",X"25",X"06",X"22",X"0A",X"A1",X"42",
		X"24",X"06",X"33",X"46",X"5A",X"26",X"F1",X"39",X"5D",X"39",X"C6",X"25",X"F7",X"A6",X"7D",X"C6",
		X"05",X"20",X"15",X"C6",X"05",X"DE",X"23",X"10",X"BE",X"BB",X"DC",X"A6",X"C4",X"A1",X"A4",X"26",
		X"07",X"AE",X"41",X"AC",X"21",X"26",X"01",X"5A",X"F7",X"A6",X"7E",X"96",X"26",X"27",X"34",X"F6",
		X"A6",X"7D",X"10",X"8E",X"A9",X"45",X"DE",X"23",X"37",X"12",X"A1",X"A4",X"26",X"20",X"AC",X"21",
		X"26",X"1C",X"7A",X"A6",X"7E",X"26",X"17",X"33",X"26",X"34",X"40",X"CC",X"AA",X"23",X"A3",X"E1",
		X"27",X"05",X"1F",X"01",X"BD",X"7F",X"33",X"7A",X"A6",X"7D",X"BD",X"E8",X"B4",X"39",X"31",X"26",
		X"5A",X"26",X"D7",X"39",X"BD",X"E0",X"EF",X"8E",X"EB",X"E2",X"BD",X"F5",X"42",X"8E",X"EC",X"05",
		X"BD",X"F5",X"42",X"86",X"B4",X"BD",X"E5",X"1F",X"4A",X"26",X"FA",X"39",X"BD",X"44",X"69",X"FD",
		X"A6",X"76",X"8E",X"E8",X"FB",X"C6",X"0E",X"8D",X"4D",X"2B",X"14",X"58",X"58",X"F7",X"A6",X"78",
		X"8E",X"E8",X"F3",X"C6",X"08",X"B6",X"A6",X"77",X"8D",X"3C",X"2B",X"03",X"FA",X"A6",X"78",X"F7",
		X"A6",X"7A",X"39",X"71",X"8B",X"8A",X"A9",X"A8",X"C7",X"C6",X"E0",X"10",X"1F",X"1E",X"30",X"2F",
		X"41",X"40",X"52",X"51",X"63",X"62",X"74",X"73",X"82",X"20",X"41",X"48",X"4F",X"56",X"42",X"49",
		X"50",X"57",X"43",X"4A",X"51",X"58",X"44",X"4B",X"52",X"59",X"45",X"4C",X"53",X"5A",X"46",X"4D",
		X"54",X"3C",X"47",X"4E",X"55",X"20",X"5A",X"2B",X"0A",X"A1",X"85",X"22",X"07",X"5A",X"A1",X"85",
		X"25",X"F4",X"54",X"39",X"5A",X"20",X"EF",X"8E",X"A6",X"51",X"EF",X"08",X"B6",X"A6",X"7B",X"2B",
		X"19",X"84",X"03",X"C6",X"1E",X"3D",X"CB",X"71",X"E7",X"02",X"B6",X"A6",X"7B",X"44",X"44",X"C6",
		X"22",X"3D",X"C3",X"00",X"20",X"ED",X"00",X"BD",X"13",X"22",X"39",X"48",X"AE",X"86",X"BD",X"F5",
		X"42",X"39",X"86",X"00",X"20",X"02",X"86",X"11",X"8E",X"A6",X"5B",X"A7",X"05",X"BD",X"F5",X"42",
		X"39",X"FE",X"A6",X"5D",X"33",X"CB",X"FF",X"A6",X"5D",X"8E",X"A6",X"62",X"6F",X"84",X"BD",X"F4",
		X"87",X"E3",X"01",X"ED",X"01",X"86",X"22",X"A7",X"84",X"BD",X"F4",X"87",X"39",X"BD",X"E9",X"62",
		X"BD",X"E9",X"9A",X"B7",X"A6",X"74",X"BD",X"E9",X"66",X"39",X"B6",X"A6",X"7B",X"8E",X"E9",X"0A",
		X"A6",X"86",X"39",X"5F",X"BD",X"E5",X"61",X"BD",X"E0",X"EC",X"4F",X"BD",X"66",X"BC",X"CC",X"0E",
		X"10",X"DD",X"55",X"8E",X"E2",X"DE",X"BF",X"AE",X"59",X"7F",X"AE",X"5B",X"8E",X"E2",X"C4",X"BF",
		X"AE",X"55",X"7F",X"AE",X"57",X"8E",X"EC",X"2D",X"BD",X"13",X"22",X"8E",X"EB",X"A7",X"BD",X"F5",
		X"4F",X"8E",X"EB",X"C6",X"BD",X"F5",X"4F",X"96",X"2C",X"27",X"08",X"8E",X"EA",X"D3",X"96",X"09",
		X"BD",X"E9",X"5B",X"4F",X"D6",X"26",X"27",X"06",X"4C",X"C1",X"25",X"2D",X"01",X"4C",X"B7",X"A6",
		X"7C",X"8E",X"EA",X"D7",X"BD",X"E9",X"5B",X"8E",X"EB",X"8D",X"BD",X"F5",X"42",X"10",X"8E",X"A6",
		X"51",X"86",X"01",X"A7",X"27",X"CC",X"01",X"03",X"ED",X"25",X"CC",X"07",X"0C",X"ED",X"23",X"8E",
		X"EC",X"21",X"AF",X"28",X"CC",X"41",X"FF",X"8E",X"A6",X"74",X"ED",X"84",X"BF",X"A6",X"5B",X"86",
		X"11",X"B7",X"A6",X"60",X"C6",X"07",X"F7",X"A6",X"79",X"C6",X"71",X"BD",X"EA",X"8E",X"C6",X"8F",
		X"BD",X"EA",X"8E",X"C6",X"AD",X"BD",X"EA",X"8E",X"C6",X"CB",X"BD",X"EA",X"8E",X"8E",X"EA",X"DD",
		X"BD",X"F5",X"4F",X"8E",X"EA",X"E7",X"BD",X"F5",X"4F",X"9E",X"23",X"86",X"03",X"5F",X"ED",X"1E",
		X"31",X"03",X"C6",X"20",X"BD",X"7F",X"26",X"CE",X"00",X"82",X"8E",X"A6",X"62",X"CC",X"22",X"58",
		X"A7",X"84",X"EF",X"01",X"E7",X"03",X"CC",X"05",X"02",X"ED",X"04",X"BD",X"F4",X"87",X"33",X"42",
		X"FF",X"A6",X"5D",X"CC",X"4D",X"20",X"B7",X"A6",X"5F",X"F7",X"A6",X"74",X"86",X"FF",X"B7",X"A6",
		X"7B",X"86",X"03",X"BD",X"E0",X"76",X"1C",X"AF",X"C6",X"08",X"BD",X"E5",X"61",X"39",X"E7",X"22",
		X"8E",X"00",X"20",X"AF",X"20",X"F6",X"A6",X"79",X"34",X"04",X"8E",X"A6",X"51",X"BD",X"13",X"22",
		X"8E",X"A6",X"5B",X"FC",X"A6",X"51",X"C3",X"00",X"09",X"ED",X"02",X"B6",X"A6",X"53",X"8B",X"07",
		X"A7",X"04",X"BD",X"F5",X"42",X"EC",X"20",X"C3",X"00",X"22",X"ED",X"20",X"B6",X"A6",X"74",X"4C",
		X"81",X"5A",X"22",X"04",X"81",X"41",X"24",X"02",X"86",X"20",X"B7",X"A6",X"74",X"6A",X"E4",X"26",
		X"C9",X"35",X"84",X"EA",X"F1",X"EB",X"00",X"EB",X"0F",X"EB",X"37",X"EB",X"60",X"EA",X"E3",X"00",
		X"D0",X"D3",X"11",X"52",X"55",X"42",X"FF",X"EA",X"ED",X"00",X"F2",X"D3",X"11",X"45",X"4E",X"44",
		X"FF",X"EA",X"F7",X"00",X"7A",X"24",X"11",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"31",X"FF",
		X"EB",X"06",X"00",X"7A",X"24",X"11",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"32",X"FF",X"EB",
		X"15",X"00",X"2F",X"31",X"22",X"59",X"4F",X"55",X"20",X"41",X"52",X"45",X"20",X"41",X"20",X"44",
		X"41",X"49",X"4C",X"59",X"20",X"54",X"55",X"52",X"4B",X"45",X"59",X"20",X"54",X"45",X"52",X"4D",
		X"49",X"4E",X"41",X"54",X"4F",X"52",X"FF",X"EB",X"3D",X"00",X"2C",X"31",X"22",X"59",X"4F",X"55",
		X"20",X"41",X"52",X"45",X"20",X"41",X"4E",X"20",X"45",X"4C",X"49",X"54",X"45",X"20",X"54",X"55",
		X"52",X"4B",X"45",X"59",X"20",X"54",X"45",X"52",X"4D",X"49",X"4E",X"41",X"54",X"4F",X"52",X"FF",
		X"EB",X"66",X"00",X"20",X"31",X"22",X"59",X"4F",X"55",X"20",X"41",X"52",X"45",X"20",X"54",X"48",
		X"45",X"20",X"47",X"52",X"45",X"41",X"54",X"45",X"53",X"54",X"20",X"54",X"55",X"52",X"4B",X"45",
		X"59",X"20",X"54",X"45",X"52",X"4D",X"49",X"4E",X"41",X"54",X"4F",X"52",X"FF",X"EB",X"93",X"00",
		X"59",X"3E",X"33",X"45",X"4E",X"54",X"45",X"52",X"20",X"59",X"4F",X"55",X"52",X"20",X"49",X"4E",
		X"49",X"54",X"49",X"41",X"4C",X"53",X"FF",X"EB",X"AD",X"00",X"22",X"62",X"44",X"41",X"49",X"4D",
		X"20",X"47",X"55",X"4E",X"20",X"54",X"4F",X"20",X"53",X"45",X"4C",X"45",X"43",X"54",X"20",X"4C",
		X"45",X"54",X"54",X"45",X"52",X"FF",X"EB",X"CC",X"00",X"A2",X"62",X"55",X"53",X"48",X"4F",X"4F",
		X"54",X"20",X"4C",X"45",X"54",X"54",X"45",X"52",X"20",X"54",X"4F",X"20",X"45",X"4E",X"54",X"45",
		X"52",X"FF",X"EB",X"E8",X"00",X"3E",X"6E",X"11",X"35",X"20",X"65",X"6E",X"74",X"72",X"69",X"65",
		X"73",X"20",X"6D",X"61",X"78",X"69",X"6D",X"75",X"6D",X"20",X"70",X"65",X"72",X"20",X"70",X"6C",
		X"61",X"79",X"65",X"72",X"FF",X"EC",X"0B",X"00",X"53",X"82",X"11",X"6C",X"6F",X"77",X"65",X"73",
		X"74",X"20",X"65",X"6E",X"74",X"72",X"79",X"20",X"72",X"65",X"70",X"6C",X"61",X"63",X"65",X"64",
		X"FF",X"EC",X"27",X"00",X"00",X"EC",X"21",X"77",X"88",X"99",X"00",X"EC",X"27",X"00",X"08",X"10",
		X"4D",X"8A",X"01",X"03",X"05",X"EC",X"37",X"EC",X"3F",X"EC",X"46",X"00",X"00",X"EC",X"37",X"BB",
		X"CC",X"DD",X"EE",X"00",X"EC",X"3F",X"EE",X"DD",X"CC",X"BB",X"00",X"EC",X"46",X"86",X"01",X"B7",
		X"C8",X"00",X"8E",X"BF",X"00",X"CC",X"2A",X"00",X"20",X"0B",X"86",X"01",X"B7",X"C8",X"00",X"8E",
		X"BB",X"B9",X"CC",X"3A",X"44",X"F7",X"C8",X"81",X"AD",X"98",X"1D",X"AD",X"98",X"1F",X"AD",X"98",
		X"21",X"86",X"06",X"B7",X"C8",X"00",X"39",X"34",X"02",X"86",X"12",X"8D",X"30",X"35",X"02",X"E6",
		X"00",X"26",X"07",X"CE",X"EC",X"F9",X"EF",X"88",X"21",X"39",X"C1",X"05",X"23",X"02",X"C6",X"05",
		X"58",X"58",X"CE",X"EC",X"BD",X"31",X"C5",X"EE",X"A1",X"EF",X"88",X"17",X"EE",X"A4",X"EF",X"88",
		X"1B",X"CE",X"EC",X"A7",X"EF",X"88",X"21",X"EE",X"88",X"17",X"FF",X"C8",X"82",X"EE",X"88",X"19",
		X"FF",X"C8",X"84",X"EE",X"88",X"1B",X"FF",X"C8",X"86",X"B7",X"C8",X"80",X"39",X"00",X"00",X"00",
		X"00",X"58",X"09",X"03",X"04",X"57",X"F1",X"03",X"08",X"57",X"CD",X"03",X"0C",X"57",X"9D",X"03",
		X"10",X"57",X"61",X"03",X"14",X"CE",X"1F",X"B7",X"FF",X"C8",X"82",X"CE",X"03",X"04",X"FF",X"C8",
		X"86",X"EE",X"88",X"13",X"FF",X"C8",X"84",X"B7",X"C8",X"80",X"39",X"34",X"02",X"86",X"12",X"8D",
		X"EA",X"CE",X"EC",X"F9",X"EF",X"88",X"1D",X"35",X"82",X"39",X"CE",X"1F",X"A3",X"FF",X"C8",X"82",
		X"CE",X"04",X"05",X"FF",X"C8",X"86",X"EE",X"88",X"15",X"FF",X"C8",X"84",X"B7",X"C8",X"80",X"39",
		X"34",X"02",X"86",X"12",X"8D",X"EA",X"CE",X"EC",X"F9",X"EF",X"88",X"1F",X"35",X"82",X"B6",X"A9",
		X"43",X"B7",X"B2",X"66",X"7F",X"B2",X"67",X"CC",X"10",X"05",X"8E",X"ED",X"FB",X"CE",X"B2",X"8A",
		X"8D",X"09",X"8E",X"EE",X"0A",X"CE",X"B2",X"FC",X"8D",X"01",X"39",X"34",X"10",X"8E",X"ED",X"F5",
		X"BD",X"F4",X"87",X"35",X"10",X"BD",X"F5",X"4F",X"8D",X"01",X"39",X"34",X"07",X"1A",X"50",X"FF",
		X"C8",X"84",X"FD",X"C8",X"86",X"7F",X"CB",X"A0",X"7F",X"C8",X"00",X"CC",X"00",X"00",X"FD",X"C8",
		X"82",X"86",X"05",X"B7",X"C8",X"80",X"CC",X"06",X"01",X"B7",X"C8",X"00",X"F7",X"CB",X"A0",X"35",
		X"87",X"DC",X"10",X"BD",X"65",X"F9",X"8E",X"B2",X"68",X"BD",X"66",X"1A",X"86",X"FF",X"A7",X"84",
		X"CC",X"06",X"05",X"8E",X"EE",X"19",X"CE",X"B2",X"6C",X"8D",X"B0",X"39",X"BD",X"65",X"F9",X"8E",
		X"B2",X"DA",X"BD",X"66",X"1A",X"86",X"FF",X"A7",X"84",X"CC",X"06",X"05",X"8E",X"EE",X"1F",X"CE",
		X"B2",X"DE",X"8D",X"97",X"39",X"B6",X"B2",X"67",X"26",X"1B",X"F6",X"A9",X"43",X"F1",X"B2",X"66",
		X"27",X"0B",X"F7",X"B2",X"66",X"8D",X"D5",X"86",X"0B",X"B7",X"B2",X"67",X"39",X"8E",X"B2",X"8A",
		X"CE",X"B2",X"6C",X"20",X"09",X"7A",X"B2",X"67",X"8E",X"B2",X"FC",X"CE",X"B2",X"DE",X"BF",X"C8",
		X"82",X"8E",X"41",X"EA",X"BF",X"C8",X"84",X"8E",X"10",X"05",X"BF",X"C8",X"86",X"86",X"06",X"B7",
		X"C8",X"80",X"8E",X"51",X"EA",X"BF",X"C8",X"84",X"8E",X"06",X"05",X"BF",X"C8",X"86",X"FF",X"C8",
		X"82",X"B7",X"C8",X"80",X"39",X"00",X"00",X"00",X"00",X"10",X"05",X"EE",X"01",X"00",X"00",X"00",
		X"BB",X"4D",X"49",X"53",X"53",X"49",X"4F",X"4E",X"20",X"FF",X"EE",X"10",X"00",X"00",X"00",X"22",
		X"43",X"52",X"45",X"44",X"49",X"54",X"53",X"20",X"FF",X"B2",X"68",X"00",X"00",X"00",X"BB",X"B2",
		X"DA",X"00",X"00",X"00",X"22",X"BD",X"E0",X"E5",X"8E",X"EE",X"DC",X"BD",X"F5",X"42",X"8D",X"5E",
		X"86",X"04",X"BD",X"E0",X"76",X"0F",X"60",X"C6",X"0A",X"CE",X"EE",X"F6",X"20",X"1C",X"B6",X"C9",
		X"80",X"85",X"01",X"27",X"15",X"86",X"EE",X"8D",X"6D",X"A6",X"04",X"5A",X"26",X"04",X"C6",X"0A",
		X"86",X"2A",X"8B",X"0C",X"A7",X"04",X"86",X"11",X"8D",X"5C",X"A6",X"C5",X"C1",X"05",X"25",X"05",
		X"BD",X"70",X"0E",X"20",X"03",X"B7",X"C9",X"86",X"86",X"1E",X"8D",X"17",X"26",X"0B",X"86",X"0C",
		X"B7",X"C9",X"86",X"86",X"1E",X"8D",X"0C",X"27",X"C5",X"CC",X"00",X"0C",X"F7",X"C9",X"86",X"BD",
		X"70",X"0E",X"39",X"BD",X"E5",X"1F",X"0D",X"60",X"26",X"03",X"4A",X"26",X"F6",X"39",X"8E",X"A8",
		X"FA",X"CC",X"00",X"7A",X"ED",X"02",X"86",X"EE",X"A7",X"05",X"CE",X"EF",X"01",X"CC",X"36",X"0A",
		X"EF",X"84",X"A7",X"04",X"BD",X"F5",X"4F",X"8B",X"0C",X"33",X"4D",X"5A",X"26",X"F2",X"CC",X"11",
		X"36",X"E7",X"04",X"8D",X"01",X"39",X"34",X"07",X"1A",X"50",X"7F",X"C8",X"00",X"B7",X"C8",X"81",
		X"86",X"3D",X"E6",X"04",X"FD",X"C8",X"82",X"FD",X"C8",X"84",X"CC",X"18",X"05",X"FD",X"C8",X"86",
		X"CC",X"06",X"1F",X"F7",X"C8",X"80",X"12",X"B7",X"C8",X"00",X"35",X"87",X"EE",X"E2",X"00",X"56",
		X"22",X"11",X"53",X"4F",X"55",X"4E",X"44",X"2D",X"43",X"4F",X"49",X"4C",X"2D",X"4C",X"41",X"4D",
		X"50",X"20",X"54",X"45",X"53",X"54",X"FF",X"1C",X"2C",X"04",X"08",X"5F",X"5E",X"5D",X"5C",X"5B",
		X"5A",X"53",X"4F",X"55",X"4E",X"44",X"20",X"4C",X"49",X"4E",X"45",X"20",X"31",X"FF",X"53",X"4F",
		X"55",X"4E",X"44",X"20",X"4C",X"49",X"4E",X"45",X"20",X"32",X"FF",X"53",X"4F",X"55",X"4E",X"44",
		X"20",X"4C",X"49",X"4E",X"45",X"20",X"33",X"FF",X"53",X"4F",X"55",X"4E",X"44",X"20",X"4C",X"49",
		X"4E",X"45",X"20",X"34",X"FF",X"53",X"4F",X"55",X"4E",X"44",X"20",X"4C",X"49",X"4E",X"45",X"20",
		X"35",X"FF",X"53",X"4F",X"55",X"4E",X"44",X"20",X"4C",X"49",X"4E",X"45",X"20",X"36",X"FF",X"47",
		X"52",X"45",X"4E",X"41",X"44",X"45",X"20",X"4C",X"41",X"4D",X"50",X"FF",X"20",X"20",X"47",X"55",
		X"4E",X"20",X"4C",X"41",X"4D",X"50",X"20",X"20",X"FF",X"46",X"45",X"41",X"54",X"48",X"45",X"52",
		X"20",X"43",X"4F",X"49",X"4C",X"FF",X"20",X"20",X"47",X"55",X"4E",X"20",X"43",X"4F",X"49",X"4C",
		X"20",X"20",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1A",X"50",X"7F",X"CB",X"80",X"7E",X"F2",X"10",X"1A",X"50",X"10",X"CE",X"BF",X"00",X"86",X"BF",
		X"1F",X"8B",X"BD",X"E0",X"E5",X"8E",X"90",X"00",X"CE",X"00",X"00",X"86",X"14",X"B7",X"C9",X"00",
		X"EF",X"81",X"8C",X"BF",X"FF",X"23",X"F6",X"BD",X"E0",X"4F",X"8E",X"10",X"80",X"CE",X"80",X"00",
		X"CC",X"03",X"10",X"B7",X"C8",X"00",X"7F",X"C8",X"81",X"BF",X"C8",X"86",X"FF",X"C8",X"84",X"F7",
		X"C8",X"80",X"86",X"06",X"B7",X"C8",X"00",X"BD",X"DB",X"0B",X"86",X"00",X"BD",X"E0",X"2D",X"BD",
		X"DF",X"C4",X"BD",X"DB",X"41",X"BD",X"F0",X"62",X"BD",X"7E",X"99",X"7E",X"D3",X"E3",X"BD",X"F0",
		X"62",X"3B",X"BD",X"DF",X"C4",X"BD",X"D1",X"41",X"BD",X"3E",X"CA",X"34",X"01",X"1A",X"50",X"4F",
		X"BD",X"66",X"BC",X"BD",X"00",X"2D",X"BD",X"E5",X"32",X"BD",X"72",X"6D",X"BD",X"14",X"01",X"BD",
		X"1B",X"51",X"7F",X"CB",X"80",X"86",X"01",X"B7",X"CB",X"A0",X"86",X"FF",X"B7",X"BC",X"2D",X"0F",
		X"E7",X"0F",X"A9",X"0F",X"9F",X"35",X"81",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",
		X"20",X"28",X"43",X"29",X"20",X"31",X"39",X"38",X"34",X"2C",X"20",X"57",X"49",X"4C",X"4C",X"49",
		X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",
		X"49",X"4E",X"43",X"2E",X"7F",X"C9",X"85",X"7F",X"C9",X"87",X"7F",X"C9",X"81",X"7F",X"C9",X"83",
		X"7F",X"C9",X"89",X"CC",X"0C",X"04",X"FD",X"C9",X"88",X"CC",X"00",X"35",X"FD",X"C9",X"84",X"CC",
		X"3C",X"05",X"FD",X"C9",X"86",X"86",X"0C",X"B7",X"C9",X"86",X"CC",X"00",X"04",X"FD",X"C9",X"80",
		X"CC",X"FF",X"3C",X"FD",X"C9",X"82",X"39",X"8E",X"F1",X"02",X"A6",X"85",X"B7",X"C9",X"8C",X"97",
		X"69",X"39",X"40",X"79",X"24",X"30",X"19",X"12",X"02",X"78",X"00",X"10",X"08",X"03",X"46",X"21",
		X"06",X"0E",X"00",X"FF",X"39",X"12",X"35",X"B2",X"35",X"CD",X"35",X"E8",X"36",X"03",X"36",X"1E",
		X"36",X"39",X"36",X"54",X"36",X"6F",X"36",X"8A",X"36",X"A5",X"36",X"C0",X"36",X"DB",X"36",X"F6",
		X"37",X"11",X"37",X"2C",X"37",X"47",X"37",X"62",X"37",X"7D",X"37",X"98",X"37",X"B3",X"37",X"CE",
		X"37",X"E9",X"38",X"04",X"38",X"1F",X"38",X"3A",X"38",X"55",X"38",X"70",X"38",X"8B",X"38",X"A6",
		X"38",X"C1",X"38",X"DC",X"38",X"F7",X"30",X"00",X"30",X"1B",X"30",X"36",X"30",X"51",X"30",X"6C",
		X"30",X"87",X"31",X"44",X"31",X"5F",X"31",X"7A",X"31",X"95",X"31",X"B0",X"31",X"CB",X"32",X"A3",
		X"32",X"BE",X"32",X"D9",X"32",X"F4",X"33",X"0F",X"33",X"CC",X"33",X"E7",X"34",X"02",X"34",X"1D",
		X"34",X"38",X"34",X"53",X"35",X"10",X"35",X"2B",X"35",X"46",X"39",X"2D",X"39",X"48",X"39",X"63",
		X"39",X"7E",X"39",X"99",X"39",X"48",X"30",X"A2",X"30",X"BD",X"30",X"D8",X"30",X"F3",X"31",X"0E",
		X"31",X"29",X"31",X"E6",X"32",X"01",X"32",X"1C",X"32",X"37",X"32",X"52",X"32",X"6D",X"33",X"45",
		X"33",X"60",X"33",X"7B",X"33",X"96",X"33",X"B1",X"34",X"6E",X"34",X"89",X"34",X"A4",X"34",X"BF",
		X"34",X"DA",X"34",X"F5",X"35",X"61",X"35",X"7C",X"35",X"97",X"BD",X"E0",X"E5",X"BD",X"E1",X"10",
		X"BD",X"D4",X"58",X"3F",X"10",X"CE",X"BF",X"00",X"8E",X"70",X"49",X"BD",X"6F",X"D3",X"B6",X"C9",
		X"80",X"85",X"01",X"26",X"1C",X"C6",X"0E",X"BD",X"E5",X"61",X"1C",X"EF",X"BD",X"FC",X"49",X"BD",
		X"FA",X"60",X"BD",X"D9",X"5E",X"BD",X"EE",X"25",X"BD",X"FD",X"58",X"BD",X"D7",X"5A",X"BD",X"D8",
		X"2D",X"BD",X"78",X"BB",X"BD",X"01",X"79",X"1A",X"50",X"10",X"CE",X"BF",X"00",X"7E",X"F0",X"08",
		X"CC",X"00",X"14",X"B7",X"C9",X"8C",X"8E",X"84",X"A8",X"F7",X"C9",X"00",X"1E",X"89",X"1E",X"89",
		X"30",X"1F",X"26",X"F5",X"86",X"06",X"B7",X"C9",X"8C",X"7F",X"C9",X"81",X"7F",X"C9",X"80",X"CE",
		X"F4",X"15",X"10",X"CE",X"F2",X"41",X"7E",X"FB",X"44",X"27",X"1B",X"7E",X"FB",X"BC",X"86",X"01",
		X"39",X"F2",X"39",X"F2",X"3E",X"F2",X"EE",X"F2",X"EE",X"F2",X"EE",X"F2",X"EE",X"F2",X"56",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"CE",X"C0",X"00",X"BD",X"F0",X"C4",X"86",X"3E",X"B7",
		X"C9",X"82",X"B6",X"C9",X"83",X"84",X"F7",X"B7",X"C9",X"83",X"8A",X"08",X"B7",X"C9",X"83",X"86",
		X"00",X"BD",X"E0",X"2D",X"86",X"38",X"BD",X"E0",X"3E",X"7F",X"C9",X"81",X"C6",X"79",X"F7",X"C9",
		X"8C",X"BD",X"FA",X"AE",X"26",X"1F",X"C6",X"24",X"F7",X"C9",X"8C",X"BD",X"FC",X"6A",X"26",X"15",
		X"86",X"40",X"B7",X"C9",X"8C",X"8E",X"F3",X"7F",X"BD",X"F5",X"42",X"8E",X"F3",X"8B",X"BD",X"F5",
		X"42",X"86",X"03",X"8D",X"10",X"C6",X"30",X"F7",X"C9",X"8C",X"BD",X"D9",X"BD",X"86",X"40",X"B7",
		X"C9",X"8C",X"7E",X"F0",X"08",X"C6",X"14",X"8E",X"84",X"A8",X"F7",X"C9",X"00",X"1E",X"89",X"1E",
		X"89",X"30",X"1F",X"26",X"F5",X"4A",X"26",X"ED",X"39",X"1A",X"50",X"10",X"CE",X"C0",X"00",X"BD",
		X"E0",X"EF",X"BD",X"FA",X"E8",X"BD",X"FA",X"D2",X"26",X"0A",X"BD",X"FC",X"79",X"26",X"05",X"BD",
		X"D9",X"70",X"27",X"F1",X"BD",X"FA",X"E8",X"10",X"CE",X"BF",X"00",X"7E",X"F0",X"08",X"7F",X"C9",
		X"81",X"CE",X"00",X"04",X"FF",X"C9",X"80",X"1F",X"43",X"10",X"CE",X"F3",X"1C",X"1F",X"02",X"7E",
		X"F3",X"32",X"1F",X"98",X"44",X"44",X"44",X"44",X"7E",X"F3",X"32",X"1F",X"98",X"84",X"0F",X"7E",
		X"F3",X"32",X"86",X"11",X"7E",X"F3",X"32",X"1F",X"20",X"1F",X"34",X"39",X"F3",X"02",X"F3",X"0B",
		X"F3",X"12",X"F3",X"17",X"34",X"01",X"1A",X"50",X"8D",X"C4",X"8D",X"C2",X"8D",X"C0",X"8D",X"BE",
		X"35",X"81",X"8E",X"F1",X"02",X"A6",X"86",X"B7",X"C9",X"8C",X"8E",X"84",X"A8",X"86",X"14",X"B7",
		X"C9",X"00",X"B6",X"C9",X"80",X"85",X"02",X"26",X"1C",X"30",X"1F",X"26",X"F0",X"86",X"FF",X"B7",
		X"C9",X"8C",X"8E",X"11",X"B0",X"86",X"14",X"B7",X"C9",X"00",X"B6",X"C9",X"80",X"85",X"02",X"26",
		X"04",X"30",X"1F",X"26",X"F0",X"39",X"86",X"05",X"B7",X"CC",X"36",X"B6",X"CC",X"36",X"84",X"0F",
		X"81",X"05",X"26",X"0A",X"73",X"CC",X"36",X"B6",X"CC",X"36",X"84",X"0F",X"81",X"0A",X"39",X"F3",
		X"91",X"00",X"4D",X"52",X"44",X"F3",X"91",X"00",X"4D",X"52",X"33",X"F3",X"A9",X"00",X"65",X"66",
		X"44",X"49",X"4E",X"49",X"54",X"49",X"41",X"4C",X"20",X"54",X"45",X"53",X"54",X"53",X"20",X"49",
		X"4E",X"44",X"49",X"43",X"41",X"54",X"45",X"3A",X"FF",X"41",X"4C",X"4C",X"20",X"53",X"59",X"53",
		X"54",X"45",X"4D",X"53",X"20",X"47",X"4F",X"21",X"FF",X"F3",X"CB",X"00",X"4A",X"78",X"11",X"F3",
		X"E4",X"00",X"56",X"87",X"11",X"F3",X"F9",X"00",X"41",X"96",X"11",X"52",X"45",X"53",X"54",X"4F",
		X"52",X"45",X"20",X"46",X"41",X"43",X"54",X"4F",X"52",X"59",X"20",X"53",X"45",X"54",X"54",X"49",
		X"4E",X"47",X"53",X"FF",X"42",X"59",X"20",X"4F",X"50",X"45",X"4E",X"49",X"4E",X"47",X"20",X"43",
		X"4F",X"49",X"4E",X"20",X"44",X"4F",X"4F",X"52",X"FF",X"41",X"4E",X"44",X"20",X"54",X"55",X"52",
		X"4E",X"49",X"4E",X"47",X"20",X"47",X"41",X"4D",X"45",X"20",X"4F",X"46",X"46",X"20",X"41",X"4E",
		X"44",X"20",X"4F",X"4E",X"FF",X"01",X"01",X"BF",X"00",X"01",X"03",X"BF",X"00",X"01",X"05",X"BF",
		X"00",X"00",X"34",X"77",X"1A",X"50",X"EC",X"81",X"FD",X"C8",X"82",X"8D",X"39",X"8D",X"4E",X"B6",
		X"BC",X"00",X"8B",X"0A",X"E6",X"61",X"F7",X"C8",X"00",X"B7",X"C8",X"80",X"C6",X"06",X"F7",X"C8",
		X"00",X"7E",X"F5",X"5E",X"34",X"77",X"1A",X"50",X"EC",X"81",X"FD",X"C8",X"82",X"8D",X"17",X"8D",
		X"2C",X"B6",X"BC",X"00",X"8B",X"0A",X"C6",X"02",X"F7",X"C8",X"00",X"B7",X"C8",X"80",X"C6",X"06",
		X"F7",X"C8",X"00",X"7E",X"F5",X"5E",X"EC",X"81",X"46",X"56",X"F7",X"C8",X"84",X"24",X"04",X"86",
		X"20",X"20",X"01",X"4F",X"B7",X"BC",X"00",X"E6",X"80",X"F7",X"C8",X"85",X"39",X"EC",X"84",X"88",
		X"00",X"C8",X"00",X"FD",X"C8",X"86",X"39",X"34",X"77",X"1A",X"50",X"A6",X"80",X"B7",X"C8",X"81",
		X"8D",X"D4",X"8D",X"E9",X"B6",X"BC",X"00",X"8B",X"12",X"B7",X"C8",X"80",X"7E",X"F5",X"5E",X"10",
		X"BF",X"BC",X"1D",X"CE",X"BC",X"01",X"ED",X"43",X"EC",X"81",X"FD",X"BC",X"21",X"EC",X"81",X"FD",
		X"BC",X"25",X"ED",X"40",X"A6",X"80",X"A7",X"42",X"A6",X"84",X"B7",X"BC",X"27",X"7F",X"BC",X"2A",
		X"7F",X"BC",X"2C",X"39",X"CE",X"BC",X"01",X"BE",X"BC",X"21",X"F6",X"BC",X"2A",X"3A",X"5C",X"F7",
		X"BC",X"2A",X"E6",X"84",X"F7",X"BC",X"2E",X"2D",X"33",X"C1",X"5C",X"26",X"0F",X"FC",X"BC",X"25",
		X"ED",X"40",X"A6",X"42",X"AB",X"44",X"8B",X"03",X"A7",X"42",X"20",X"25",X"8D",X"24",X"EC",X"40",
		X"FD",X"BC",X"2F",X"A6",X"42",X"B7",X"BC",X"31",X"1F",X"31",X"BD",X"F4",X"66",X"BD",X"F4",X"7D",
		X"8D",X"22",X"4F",X"E6",X"43",X"58",X"E3",X"40",X"ED",X"40",X"20",X"05",X"86",X"FF",X"B7",X"BC",
		X"2C",X"39",X"BE",X"BC",X"1D",X"C0",X"20",X"58",X"3A",X"AE",X"84",X"BF",X"C8",X"82",X"39",X"BE",
		X"BC",X"1F",X"20",X"F1",X"B6",X"BC",X"28",X"B7",X"C8",X"81",X"B6",X"BC",X"00",X"8B",X"1A",X"C6",
		X"02",X"F7",X"C8",X"00",X"B7",X"C8",X"80",X"C6",X"06",X"F7",X"C8",X"00",X"39",X"B6",X"BC",X"29",
		X"20",X"E5",X"34",X"77",X"1A",X"50",X"CC",X"03",X"09",X"10",X"8E",X"F1",X"14",X"20",X"0B",X"34",
		X"77",X"1A",X"50",X"CC",X"02",X"05",X"10",X"8E",X"0A",X"33",X"8D",X"04",X"8D",X"21",X"35",X"F7",
		X"10",X"BF",X"BC",X"1F",X"CE",X"BC",X"06",X"ED",X"43",X"EC",X"81",X"FD",X"BC",X"23",X"EC",X"81",
		X"ED",X"40",X"A6",X"80",X"A7",X"42",X"A6",X"84",X"B7",X"BC",X"29",X"7F",X"BC",X"2B",X"39",X"BE",
		X"BC",X"23",X"F6",X"BC",X"2B",X"3A",X"5C",X"F7",X"BC",X"2B",X"E6",X"84",X"2D",X"18",X"BD",X"F5",
		X"1F",X"1F",X"31",X"BD",X"F4",X"66",X"BD",X"F4",X"7D",X"BD",X"F5",X"3D",X"4F",X"E6",X"43",X"58",
		X"E3",X"40",X"ED",X"40",X"20",X"D9",X"39",X"34",X"77",X"1A",X"50",X"1F",X"13",X"10",X"8E",X"BC",
		X"32",X"8E",X"00",X"96",X"86",X"05",X"BD",X"DF",X"A0",X"FC",X"BC",X"32",X"A3",X"63",X"C3",X"BC",
		X"32",X"FD",X"BC",X"32",X"8E",X"BC",X"32",X"BD",X"F5",X"CC",X"35",X"F7",X"34",X"77",X"1A",X"50",
		X"CC",X"03",X"01",X"D7",X"F1",X"B7",X"BC",X"2D",X"CE",X"BC",X"10",X"6F",X"40",X"CC",X"03",X"09",
		X"ED",X"44",X"CE",X"BC",X"0B",X"ED",X"43",X"CE",X"BC",X"16",X"ED",X"45",X"CC",X"3C",X"75",X"ED",
		X"40",X"10",X"8E",X"F1",X"14",X"CC",X"03",X"09",X"BD",X"F4",X"9F",X"35",X"F7",X"B6",X"BC",X"2D",
		X"2D",X"20",X"0A",X"F1",X"26",X"0A",X"86",X"04",X"97",X"F1",X"8E",X"70",X"D9",X"BD",X"6F",X"D3",
		X"B6",X"BC",X"2D",X"4C",X"81",X"01",X"23",X"01",X"4F",X"B7",X"BC",X"2D",X"48",X"8E",X"F6",X"23",
		X"AD",X"96",X"39",X"F6",X"27",X"F6",X"55",X"8D",X"03",X"8D",X"19",X"39",X"96",X"29",X"81",X"02",
		X"27",X"11",X"CE",X"BC",X"01",X"8E",X"BC",X"10",X"EC",X"40",X"ED",X"01",X"A6",X"42",X"A7",X"03",
		X"BD",X"F4",X"87",X"39",X"86",X"DD",X"B7",X"BC",X"28",X"BD",X"F4",X"C4",X"B6",X"BC",X"2C",X"27",
		X"03",X"B7",X"BC",X"2D",X"39",X"8D",X"03",X"8D",X"19",X"39",X"96",X"29",X"81",X"02",X"27",X"11",
		X"CE",X"BC",X"01",X"8E",X"BC",X"16",X"EC",X"40",X"ED",X"02",X"A6",X"42",X"A7",X"04",X"BD",X"F4",
		X"44",X"39",X"F6",X"BC",X"2E",X"C1",X"5C",X"27",X"1F",X"BD",X"F5",X"12",X"8E",X"BC",X"0B",X"FC",
		X"BC",X"2F",X"ED",X"00",X"B6",X"BC",X"31",X"A7",X"02",X"BD",X"F4",X"66",X"BD",X"F4",X"7D",X"B6",
		X"BC",X"27",X"B7",X"BC",X"28",X"BD",X"F5",X"24",X"39",X"CE",X"90",X"00",X"BD",X"F6",X"E5",X"FF",
		X"BB",X"97",X"39",X"FE",X"BB",X"97",X"27",X"03",X"BD",X"F7",X"29",X"39",X"CE",X"90",X"60",X"BD",
		X"F6",X"E5",X"FF",X"BB",X"93",X"39",X"FE",X"BB",X"93",X"27",X"03",X"BD",X"F7",X"29",X"39",X"CE",
		X"90",X"00",X"BD",X"F8",X"48",X"FF",X"BB",X"99",X"39",X"FE",X"BB",X"99",X"27",X"03",X"BD",X"F8",
		X"80",X"39",X"CE",X"90",X"60",X"BD",X"F8",X"48",X"FF",X"BB",X"95",X"39",X"FE",X"BB",X"95",X"27",
		X"03",X"BD",X"F8",X"80",X"39",X"4F",X"B7",X"C8",X"81",X"A7",X"45",X"D6",X"29",X"C1",X"02",X"10",
		X"27",X"00",X"C8",X"97",X"5E",X"EE",X"C8",X"12",X"27",X"2E",X"EC",X"44",X"C1",X"80",X"24",X"28",
		X"FD",X"C8",X"84",X"AE",X"46",X"BF",X"C8",X"86",X"AD",X"D8",X"0A",X"A6",X"4F",X"27",X"07",X"86",
		X"12",X"B7",X"C8",X"80",X"6F",X"4F",X"A6",X"45",X"A0",X"C8",X"2A",X"91",X"5E",X"24",X"D4",X"D6",
		X"5D",X"26",X"D0",X"BD",X"F7",X"73",X"26",X"D2",X"39",X"7F",X"C8",X"81",X"D6",X"29",X"C1",X"02",
		X"10",X"27",X"00",X"D5",X"AE",X"C8",X"10",X"A6",X"05",X"AB",X"88",X"2A",X"97",X"5E",X"20",X"08",
		X"97",X"5E",X"EE",X"C8",X"12",X"26",X"01",X"39",X"AE",X"44",X"BF",X"C8",X"84",X"AE",X"46",X"BF",
		X"C8",X"86",X"AD",X"D8",X"0A",X"A6",X"4F",X"27",X"07",X"86",X"12",X"B7",X"C8",X"80",X"6F",X"4F",
		X"A6",X"45",X"A0",X"C8",X"2A",X"91",X"5E",X"24",X"D7",X"D6",X"5D",X"26",X"D3",X"BD",X"F7",X"73",
		X"26",X"D6",X"39",X"AE",X"C8",X"10",X"0C",X"5D",X"A6",X"45",X"A0",X"C8",X"2A",X"1F",X"89",X"10",
		X"AE",X"C8",X"12",X"10",X"AF",X"88",X"12",X"10",X"BF",X"BB",X"91",X"26",X"04",X"10",X"AE",X"C8",
		X"20",X"AF",X"A8",X"10",X"AE",X"88",X"10",X"1F",X"98",X"A0",X"05",X"AB",X"88",X"2A",X"25",X"F4",
		X"10",X"AE",X"88",X"12",X"EF",X"88",X"12",X"AF",X"C8",X"10",X"10",X"AF",X"C8",X"12",X"26",X"04",
		X"10",X"AE",X"C8",X"20",X"EF",X"A8",X"10",X"FE",X"BB",X"91",X"39",X"EE",X"C8",X"12",X"27",X"42",
		X"EC",X"44",X"C1",X"80",X"24",X"3C",X"FD",X"C8",X"84",X"AE",X"42",X"BF",X"C8",X"82",X"A6",X"C8",
		X"1F",X"AE",X"46",X"BF",X"C8",X"86",X"E6",X"40",X"34",X"06",X"86",X"06",X"B7",X"C8",X"00",X"AD",
		X"D8",X"0A",X"35",X"06",X"6D",X"4F",X"27",X"0C",X"B7",X"C8",X"00",X"C4",X"20",X"CA",X"1A",X"F7",
		X"C8",X"80",X"6F",X"4F",X"A6",X"45",X"AE",X"C8",X"10",X"A1",X"05",X"24",X"BE",X"BD",X"F7",X"78",
		X"26",X"BE",X"39",X"EE",X"C8",X"12",X"26",X"01",X"39",X"AE",X"42",X"BF",X"C8",X"82",X"A6",X"C8",
		X"1F",X"AE",X"44",X"BF",X"C8",X"84",X"AE",X"46",X"BF",X"C8",X"86",X"E6",X"40",X"34",X"06",X"86",
		X"06",X"B7",X"C8",X"00",X"AD",X"D8",X"0A",X"35",X"06",X"6D",X"4F",X"27",X"0C",X"B7",X"C8",X"00",
		X"C4",X"20",X"CA",X"1A",X"F7",X"C8",X"80",X"6F",X"4F",X"A6",X"45",X"AE",X"C8",X"10",X"A1",X"05",
		X"24",X"C1",X"BD",X"F7",X"78",X"26",X"C2",X"39",X"34",X"19",X"EE",X"C8",X"12",X"27",X"2F",X"10",
		X"FF",X"BB",X"9D",X"7A",X"C9",X"85",X"7A",X"C9",X"87",X"A6",X"45",X"81",X"62",X"22",X"0E",X"A6",
		X"C8",X"1F",X"B7",X"C8",X"00",X"37",X"7F",X"34",X"3F",X"EE",X"48",X"26",X"EC",X"10",X"FE",X"BB",
		X"9D",X"86",X"06",X"B7",X"C8",X"00",X"1A",X"50",X"7C",X"C9",X"85",X"7C",X"C9",X"87",X"35",X"99",
		X"34",X"59",X"10",X"FF",X"BB",X"9D",X"7A",X"C9",X"85",X"7A",X"C9",X"87",X"A6",X"C8",X"1F",X"B7",
		X"C8",X"00",X"37",X"7F",X"34",X"3F",X"EE",X"48",X"26",X"F2",X"1A",X"50",X"7C",X"C9",X"85",X"7C",
		X"C9",X"87",X"86",X"06",X"B7",X"C8",X"00",X"10",X"FE",X"BB",X"9D",X"35",X"D9",X"34",X"37",X"10",
		X"8E",X"F8",X"F2",X"20",X"06",X"34",X"37",X"10",X"8E",X"F8",X"F8",X"BE",X"BA",X"1D",X"EE",X"81",
		X"27",X"2A",X"BF",X"BA",X"1D",X"BE",X"BA",X"9D",X"EF",X"83",X"BF",X"BA",X"9D",X"EC",X"A4",X"A7",
		X"4E",X"E7",X"C8",X"24",X"AE",X"22",X"AF",X"C8",X"20",X"AE",X"24",X"AF",X"C8",X"22",X"35",X"01",
		X"4F",X"A7",X"4C",X"A7",X"4F",X"A7",X"C8",X"2A",X"A7",X"41",X"35",X"B6",X"35",X"01",X"86",X"FF",
		X"35",X"B6",X"01",X"00",X"90",X"00",X"F9",X"12",X"01",X"02",X"90",X"60",X"F9",X"16",X"34",X"41",
		X"1A",X"50",X"8D",X"A9",X"20",X"06",X"34",X"41",X"1A",X"50",X"8D",X"A9",X"A7",X"4C",X"8D",X"23",
		X"35",X"C1",X"34",X"11",X"20",X"02",X"34",X"11",X"1A",X"50",X"6D",X"C8",X"24",X"2B",X"0F",X"BE",
		X"BB",X"1D",X"EF",X"83",X"BF",X"BB",X"1D",X"8D",X"07",X"86",X"FF",X"A7",X"C8",X"24",X"35",X"91",
		X"8E",X"F9",X"CA",X"AF",X"4A",X"CC",X"12",X"00",X"ED",X"40",X"8E",X"01",X"01",X"AF",X"46",X"CC",
		X"01",X"05",X"ED",X"4E",X"E7",X"C8",X"1F",X"6F",X"C8",X"1D",X"39",X"34",X"10",X"6D",X"C8",X"24",
		X"2B",X"05",X"AE",X"C8",X"22",X"AF",X"4A",X"35",X"90",X"96",X"40",X"26",X"6E",X"BE",X"BA",X"9D",
		X"10",X"AE",X"81",X"27",X"65",X"BF",X"BA",X"9D",X"EE",X"A8",X"20",X"4F",X"A7",X"2F",X"A7",X"45",
		X"A6",X"25",X"81",X"80",X"24",X"32",X"EE",X"C8",X"12",X"26",X"16",X"EF",X"A8",X"12",X"EE",X"A8",
		X"20",X"AE",X"C8",X"10",X"AF",X"A8",X"10",X"10",X"AF",X"C8",X"10",X"10",X"AF",X"88",X"12",X"20",
		X"34",X"A1",X"45",X"22",X"E1",X"EF",X"A8",X"12",X"AE",X"C8",X"10",X"AF",X"A8",X"10",X"10",X"AF",
		X"C8",X"10",X"10",X"AF",X"88",X"12",X"20",X"1D",X"EE",X"C8",X"10",X"A1",X"45",X"25",X"F9",X"AE",
		X"C8",X"12",X"EF",X"A8",X"10",X"10",X"AF",X"C8",X"12",X"AF",X"A8",X"12",X"26",X"03",X"AE",X"A8",
		X"20",X"10",X"AF",X"88",X"10",X"BD",X"7D",X"F5",X"86",X"FF",X"39",X"4F",X"39",X"BE",X"BB",X"1D",
		X"EE",X"81",X"27",X"21",X"BF",X"BB",X"1D",X"AE",X"C8",X"12",X"10",X"AE",X"C8",X"10",X"AF",X"A8",
		X"12",X"26",X"03",X"AE",X"C8",X"20",X"10",X"AF",X"88",X"10",X"BE",X"BA",X"1D",X"EF",X"83",X"BF",
		X"BA",X"1D",X"BD",X"7E",X"1B",X"39",X"34",X"36",X"BE",X"BA",X"9D",X"10",X"BE",X"BA",X"1D",X"20",
		X"05",X"BF",X"BA",X"9D",X"ED",X"A3",X"EC",X"81",X"26",X"F7",X"10",X"BF",X"BA",X"1D",X"35",X"B6",
		X"CE",X"90",X"00",X"8E",X"00",X"00",X"EF",X"C8",X"10",X"AF",X"C8",X"12",X"BF",X"BB",X"97",X"BF",
		X"BB",X"99",X"CE",X"90",X"60",X"EF",X"C8",X"10",X"AF",X"C8",X"12",X"BF",X"BB",X"93",X"BF",X"BB",
		X"95",X"CE",X"BA",X"1F",X"EF",X"5E",X"8E",X"90",X"C0",X"86",X"38",X"10",X"8E",X"C8",X"88",X"10",
		X"AF",X"08",X"AF",X"C1",X"30",X"88",X"60",X"4A",X"26",X"F1",X"CC",X"00",X"00",X"ED",X"C4",X"CE",
		X"BB",X"0F",X"ED",X"C4",X"FF",X"BA",X"9D",X"CE",X"BB",X"8F",X"ED",X"C4",X"FF",X"BB",X"1D",X"39",
		X"1A",X"50",X"35",X"40",X"DF",X"00",X"10",X"CE",X"C0",X"00",X"BD",X"E0",X"EF",X"BD",X"FA",X"E8",
		X"BD",X"FA",X"FE",X"26",X"1E",X"BD",X"FB",X"21",X"26",X"19",X"BD",X"FB",X"2F",X"26",X"14",X"B6",
		X"C9",X"80",X"85",X"02",X"27",X"EA",X"BD",X"FB",X"F2",X"8E",X"FC",X"11",X"BD",X"F5",X"42",X"8D",
		X"3B",X"20",X"02",X"8D",X"34",X"10",X"CE",X"BF",X"00",X"3F",X"0F",X"60",X"C6",X"0E",X"BD",X"E5",
		X"61",X"1C",X"EF",X"BD",X"E5",X"1F",X"0D",X"60",X"27",X"F9",X"DE",X"00",X"6E",X"C4",X"1A",X"50",
		X"BD",X"FA",X"FE",X"26",X"14",X"BD",X"E1",X"10",X"BD",X"FB",X"21",X"26",X"0C",X"BD",X"FB",X"2F",
		X"26",X"07",X"BD",X"E0",X"EF",X"8D",X"05",X"4F",X"39",X"BD",X"FB",X"D7",X"86",X"06",X"B7",X"C8",
		X"00",X"39",X"BD",X"FA",X"FE",X"26",X"0E",X"BD",X"FB",X"21",X"26",X"09",X"BD",X"FB",X"2F",X"26",
		X"04",X"8D",X"E9",X"4F",X"39",X"8D",X"E2",X"39",X"7F",X"C9",X"81",X"CC",X"00",X"04",X"FD",X"C9",
		X"80",X"C6",X"14",X"B6",X"C9",X"80",X"F7",X"C9",X"00",X"85",X"02",X"26",X"F6",X"39",X"CE",X"FC",
		X"2E",X"86",X"03",X"B7",X"C8",X"00",X"8D",X"3C",X"27",X"16",X"E8",X"A4",X"86",X"61",X"C5",X"F0",
		X"26",X"01",X"4C",X"1E",X"20",X"C5",X"01",X"1E",X"20",X"27",X"02",X"8B",X"02",X"1F",X"89",X"5D",
		X"39",X"CE",X"FC",X"33",X"7F",X"C8",X"00",X"BD",X"FB",X"44",X"27",X"02",X"C6",X"43",X"39",X"CE",
		X"FC",X"38",X"86",X"06",X"BD",X"E0",X"76",X"7F",X"C8",X"00",X"BD",X"FB",X"44",X"27",X"04",X"BD",
		X"FB",X"BC",X"5D",X"39",X"37",X"26",X"4D",X"27",X"60",X"1F",X"8B",X"4F",X"8E",X"01",X"00",X"58",
		X"46",X"24",X"04",X"88",X"1D",X"C8",X"87",X"ED",X"A1",X"30",X"1E",X"26",X"F2",X"1F",X"01",X"86",
		X"14",X"B7",X"C9",X"00",X"B6",X"C9",X"80",X"85",X"02",X"26",X"3E",X"1F",X"B8",X"4A",X"1F",X"8B",
		X"1F",X"10",X"26",X"D8",X"10",X"AE",X"5E",X"EC",X"5C",X"1F",X"8B",X"4F",X"8E",X"01",X"00",X"58",
		X"46",X"24",X"04",X"88",X"1D",X"C8",X"87",X"10",X"A3",X"A1",X"26",X"23",X"30",X"1E",X"26",X"EF",
		X"1F",X"01",X"86",X"14",X"B7",X"C9",X"00",X"B6",X"C9",X"80",X"85",X"02",X"26",X"0B",X"1F",X"B8",
		X"4A",X"1F",X"8B",X"1F",X"10",X"26",X"D5",X"20",X"9B",X"86",X"BF",X"1F",X"8B",X"4F",X"39",X"E1",
		X"A2",X"26",X"04",X"1F",X"89",X"E1",X"A2",X"86",X"BF",X"1F",X"8B",X"39",X"E8",X"A4",X"4F",X"1E",
		X"20",X"80",X"03",X"24",X"FC",X"8B",X"04",X"5F",X"31",X"AB",X"1E",X"20",X"48",X"48",X"48",X"48",
		X"4C",X"56",X"24",X"FC",X"1F",X"89",X"39",X"34",X"04",X"8D",X"17",X"A6",X"E4",X"C6",X"AA",X"8E",
		X"FC",X"01",X"BD",X"FC",X"A0",X"35",X"04",X"86",X"01",X"BD",X"F3",X"24",X"86",X"06",X"B7",X"C8",
		X"00",X"39",X"34",X"06",X"BD",X"E0",X"EF",X"BD",X"E1",X"10",X"86",X"04",X"BD",X"E0",X"76",X"35",
		X"86",X"FC",X"07",X"00",X"6E",X"66",X"33",X"52",X"41",X"4D",X"20",X"45",X"52",X"52",X"4F",X"52",
		X"FF",X"FC",X"17",X"00",X"50",X"66",X"44",X"4E",X"4F",X"20",X"52",X"41",X"4D",X"20",X"45",X"52",
		X"52",X"4F",X"52",X"53",X"20",X"44",X"45",X"54",X"45",X"43",X"54",X"45",X"44",X"FF",X"08",X"15",
		X"80",X"00",X"00",X"08",X"15",X"C0",X"00",X"00",X"BF",X"FF",X"00",X"00",X"BF",X"F8",X"00",X"00",
		X"BF",X"FE",X"00",X"00",X"BF",X"FC",X"00",X"00",X"00",X"0F",X"60",X"8D",X"34",X"27",X"0C",X"BD",
		X"FC",X"8D",X"1F",X"89",X"86",X"02",X"BD",X"F3",X"24",X"20",X"07",X"8E",X"FD",X"3B",X"BD",X"F5",
		X"42",X"5F",X"BD",X"E5",X"1F",X"0D",X"60",X"27",X"F9",X"39",X"BD",X"FC",X"81",X"27",X"09",X"8D",
		X"1C",X"1F",X"89",X"86",X"02",X"BD",X"F3",X"24",X"39",X"8D",X"EF",X"27",X"03",X"BD",X"F3",X"24",
		X"39",X"BD",X"E0",X"EF",X"86",X"04",X"BD",X"E0",X"76",X"BD",X"FC",X"EC",X"39",X"C6",X"F0",X"CB",
		X"10",X"80",X"0A",X"24",X"FA",X"8B",X"0A",X"34",X"04",X"AA",X"E0",X"8E",X"FD",X"2B",X"C6",X"AA",
		X"34",X"16",X"BD",X"E0",X"E5",X"BD",X"E1",X"10",X"86",X"04",X"BD",X"E0",X"76",X"B6",X"C9",X"81",
		X"85",X"04",X"26",X"06",X"8E",X"F3",X"85",X"BD",X"F5",X"42",X"35",X"16",X"BD",X"F5",X"42",X"34",
		X"02",X"32",X"77",X"30",X"63",X"10",X"EF",X"84",X"6F",X"02",X"E7",X"03",X"C6",X"66",X"E7",X"04",
		X"C6",X"33",X"E7",X"05",X"1F",X"89",X"44",X"44",X"44",X"44",X"C4",X"0F",X"C3",X"30",X"30",X"ED",
		X"1D",X"86",X"FF",X"A7",X"1F",X"BD",X"F5",X"42",X"32",X"69",X"35",X"82",X"34",X"01",X"1A",X"50",
		X"10",X"8E",X"FF",X"BA",X"8E",X"3E",X"E4",X"5F",X"20",X"09",X"A6",X"A0",X"27",X"29",X"84",X"E0",
		X"5F",X"1F",X"01",X"A6",X"A0",X"B7",X"C8",X"00",X"84",X"F8",X"1F",X"03",X"5C",X"E9",X"C0",X"30",
		X"1C",X"26",X"FA",X"BD",X"DF",X"C4",X"E1",X"A0",X"27",X"E0",X"A6",X"3D",X"84",X"1F",X"C6",X"06",
		X"F7",X"C8",X"00",X"35",X"01",X"5D",X"39",X"35",X"01",X"5F",X"39",X"FD",X"31",X"00",X"6E",X"66",
		X"33",X"52",X"4F",X"4D",X"20",X"45",X"52",X"52",X"4F",X"52",X"FF",X"FD",X"41",X"00",X"50",X"66",
		X"44",X"4E",X"4F",X"20",X"52",X"4F",X"4D",X"20",X"45",X"52",X"52",X"4F",X"52",X"53",X"20",X"44",
		X"45",X"54",X"45",X"43",X"54",X"45",X"44",X"FF",X"BD",X"E0",X"E5",X"8E",X"FF",X"0D",X"BD",X"F5",
		X"42",X"8E",X"FE",X"C1",X"BD",X"F5",X"4F",X"8E",X"FE",X"E8",X"BD",X"F5",X"4F",X"8D",X"22",X"86",
		X"04",X"BD",X"E0",X"76",X"86",X"3C",X"97",X"B5",X"BD",X"E5",X"1F",X"8D",X"14",X"B6",X"C9",X"80",
		X"85",X"02",X"27",X"F0",X"96",X"B5",X"26",X"F0",X"39",X"CB",X"09",X"F1",X"CB",X"E0",X"22",X"FB",
		X"39",X"7F",X"BB",X"E3",X"CE",X"FE",X"97",X"10",X"8E",X"BB",X"E7",X"86",X"1D",X"B7",X"BB",X"E5",
		X"F6",X"C9",X"80",X"8D",X"24",X"F6",X"C9",X"86",X"8D",X"1F",X"F6",X"C9",X"84",X"C4",X"80",X"C8",
		X"80",X"BD",X"F3",X"66",X"27",X"02",X"CA",X"01",X"8D",X"0F",X"86",X"35",X"8E",X"FE",X"F7",X"8D",
		X"44",X"86",X"3D",X"8E",X"FE",X"D2",X"8D",X"3D",X"39",X"34",X"04",X"A6",X"C0",X"27",X"34",X"C6",
		X"EE",X"A4",X"E4",X"27",X"0C",X"C6",X"11",X"A1",X"A4",X"27",X"06",X"8E",X"70",X"DD",X"BD",X"6F",
		X"D3",X"A7",X"A0",X"B6",X"BB",X"E5",X"8B",X"0B",X"FD",X"BB",X"E5",X"AE",X"C1",X"BF",X"BB",X"E1",
		X"C6",X"94",X"C0",X"02",X"6D",X"80",X"2A",X"FA",X"F7",X"BB",X"E4",X"8E",X"BB",X"E1",X"BD",X"F5",
		X"4F",X"20",X"C8",X"35",X"84",X"34",X"01",X"1A",X"50",X"B7",X"C9",X"85",X"B6",X"C9",X"84",X"35",
		X"01",X"C6",X"06",X"34",X"06",X"48",X"48",X"EE",X"06",X"C6",X"30",X"48",X"24",X"02",X"C6",X"31",
		X"E7",X"C0",X"6A",X"61",X"26",X"F3",X"C6",X"FF",X"E7",X"C0",X"E6",X"03",X"BD",X"FD",X"89",X"BD",
		X"F4",X"87",X"30",X"06",X"BD",X"F5",X"42",X"30",X"06",X"34",X"01",X"1A",X"50",X"EE",X"00",X"FF",
		X"C8",X"82",X"EE",X"02",X"FF",X"C8",X"86",X"CC",X"DD",X"05",X"B7",X"C8",X"81",X"CE",X"47",X"0D",
		X"A6",X"61",X"84",X"3F",X"A6",X"C6",X"F7",X"C8",X"00",X"E6",X"08",X"EE",X"04",X"A7",X"61",X"27",
		X"02",X"8D",X"14",X"86",X"AA",X"B7",X"C8",X"81",X"86",X"3F",X"A0",X"61",X"27",X"02",X"8D",X"07",
		X"86",X"06",X"B7",X"C8",X"00",X"35",X"87",X"34",X"02",X"86",X"1A",X"EB",X"09",X"F7",X"C8",X"85",
		X"1E",X"03",X"E3",X"06",X"B7",X"C8",X"84",X"5D",X"1E",X"03",X"2A",X"02",X"8A",X"20",X"B7",X"C8",
		X"80",X"6A",X"E4",X"26",X"E4",X"35",X"82",X"02",X"FF",X"1F",X"01",X"FF",X"27",X"04",X"FF",X"2F",
		X"08",X"FF",X"3E",X"10",X"FF",X"48",X"20",X"FF",X"54",X"40",X"FF",X"5F",X"00",X"40",X"FF",X"69",
		X"80",X"FF",X"78",X"02",X"FF",X"87",X"01",X"FF",X"8E",X"00",X"80",X"FF",X"96",X"01",X"FF",X"9B",
		X"00",X"FE",X"C7",X"00",X"7E",X"C1",X"11",X"48",X"4F",X"52",X"49",X"5A",X"4F",X"4E",X"54",X"41",
		X"4C",X"FF",X"00",X"00",X"80",X"CA",X"12",X"07",X"BB",X"F4",X"00",X"80",X"CA",X"11",X"58",X"32",
		X"02",X"10",X"19",X"00",X"01",X"80",X"D6",X"00",X"FE",X"EE",X"00",X"28",X"74",X"11",X"56",X"45",
		X"52",X"54",X"49",X"43",X"41",X"4C",X"FF",X"00",X"00",X"26",X"7D",X"12",X"07",X"BB",X"F4",X"00",
		X"26",X"7D",X"11",X"58",X"22",X"08",X"02",X"0A",X"00",X"00",X"00",X"1D",X"03",X"FF",X"13",X"00",
		X"71",X"16",X"11",X"53",X"57",X"49",X"54",X"43",X"48",X"20",X"54",X"45",X"53",X"54",X"FF",X"41",
		X"44",X"56",X"41",X"4E",X"43",X"45",X"FF",X"41",X"55",X"54",X"4F",X"20",X"55",X"50",X"FF",X"48",
		X"49",X"2D",X"53",X"43",X"4F",X"52",X"45",X"20",X"52",X"45",X"53",X"45",X"54",X"FF",X"4C",X"45",
		X"46",X"54",X"20",X"43",X"4F",X"49",X"4E",X"FF",X"43",X"45",X"4E",X"54",X"45",X"52",X"20",X"43",
		X"4F",X"49",X"4E",X"FF",X"52",X"49",X"47",X"48",X"54",X"20",X"43",X"4F",X"49",X"4E",X"FF",X"53",
		X"4C",X"41",X"4D",X"2F",X"54",X"49",X"4C",X"54",X"FF",X"31",X"20",X"50",X"4C",X"41",X"59",X"45",
		X"52",X"20",X"53",X"54",X"41",X"52",X"54",X"FF",X"32",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",
		X"20",X"53",X"54",X"41",X"52",X"54",X"FF",X"47",X"4F",X"42",X"42",X"4C",X"45",X"FF",X"47",X"52",
		X"45",X"4E",X"41",X"44",X"45",X"FF",X"46",X"49",X"52",X"45",X"FF",X"43",X"4F",X"49",X"4E",X"20",
		X"44",X"4F",X"4F",X"52",X"20",X"43",X"4C",X"4F",X"53",X"45",X"44",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"43",X"F6",X"5E",X"8B",X"01",X"B2",X"89",
		X"21",X"B3",X"87",X"41",X"33",X"85",X"61",X"54",X"91",X"02",X"94",X"8F",X"22",X"D6",X"8A",X"05",
		X"EC",X"88",X"25",X"65",X"86",X"45",X"D3",X"84",X"65",X"F1",X"42",X"E6",X"4A",X"32",X"DE",X"43",
		X"32",X"D6",X"80",X"90",X"06",X"12",X"8E",X"26",X"C8",X"8D",X"46",X"36",X"8C",X"66",X"A1",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E4",X"80",X"E4",X"3C",X"F0",X"5E",X"00",X"00",X"F0",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
