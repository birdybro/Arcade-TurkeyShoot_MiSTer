library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity turkey_shoot_bank_d is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of turkey_shoot_bank_d is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"DC",X"C0",X"0C",X"00",X"00",X"00",X"DC",X"CF",X"CC",X"FC",X"CC",X"00",X"00",
		X"00",X"0D",X"CC",X"CC",X"CC",X"D0",X"00",X"00",X"00",X"00",X"CD",X"DC",X"CC",X"CD",X"00",X"00",
		X"00",X"00",X"DC",X"FF",X"FC",X"CD",X"00",X"00",X"00",X"0C",X"CD",X"CF",X"FD",X"C0",X"00",X"00",
		X"00",X"CC",X"CC",X"CC",X"CC",X"CC",X"00",X"00",X"00",X"D0",X"0C",X"DC",X"CF",X"CC",X"C0",X"00",
		X"00",X"00",X"CC",X"CD",X"DF",X"FC",X"00",X"00",X"00",X"00",X"CC",X"0C",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"DD",X"00",X"00",X"CD",X"00",X"00",X"00",X"00",
		X"CC",X"00",X"D0",X"00",X"0D",X"0C",X"C0",X"00",X"0C",X"00",X"09",X"9A",X"A0",X"0C",X"00",X"00",
		X"00",X"0C",X"CE",X"FF",X"DA",X"00",X"00",X"00",X"00",X"0C",X"CF",X"CC",X"CF",X"CC",X"0D",X"00",
		X"00",X"09",X"EF",X"CC",X"CF",X"CC",X"00",X"00",X"0C",X"C9",X"CF",X"FF",X"FF",X"DD",X"00",X"00",
		X"DC",X"CD",X"CF",X"CC",X"FF",X"A0",X"0C",X"00",X"0D",X"00",X"DE",X"CC",X"FC",X"C0",X"00",X"00",
		X"00",X"00",X"09",X"9A",X"A0",X"C0",X"00",X"00",X"00",X"0C",X"C0",X"00",X"00",X"00",X"C0",X"00",
		X"00",X"0D",X"C0",X"00",X"D0",X"0C",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"9A",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"9E",X"FF",X"FA",X"00",X"00",X"00",X"00",X"09",X"EF",X"FF",X"FF",X"A0",X"00",X"00",
		X"00",X"09",X"EF",X"FF",X"FF",X"A0",X"00",X"00",X"00",X"09",X"4F",X"FF",X"FF",X"A0",X"00",X"00",
		X"00",X"09",X"EF",X"FF",X"FF",X"A0",X"00",X"00",X"00",X"00",X"9E",X"FF",X"FA",X"00",X"00",X"00",
		X"00",X"00",X"09",X"9A",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"66",X"66",X"66",X"66",X"00",X"00",X"06",X"67",
		X"73",X"36",X"66",X"60",X"00",X"06",X"77",X"33",X"33",X"66",X"60",X"00",X"66",X"73",X"33",X"36",
		X"66",X"66",X"00",X"63",X"33",X"66",X"66",X"66",X"66",X"00",X"63",X"33",X"36",X"66",X"66",X"66",
		X"00",X"63",X"33",X"33",X"66",X"66",X"66",X"00",X"03",X"33",X"33",X"33",X"66",X"60",X"00",X"03",
		X"33",X"33",X"33",X"66",X"60",X"00",X"00",X"33",X"32",X"26",X"66",X"00",X"00",X"00",X"00",X"66",
		X"66",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"00",X"00",X"00",X"00",X"55",X"55",X"55",X"55",
		X"00",X"00",X"05",X"50",X"04",X"45",X"55",X"50",X"00",X"05",X"00",X"44",X"45",X"55",X"50",X"00",
		X"55",X"04",X"44",X"45",X"55",X"55",X"00",X"54",X"44",X"55",X"55",X"55",X"55",X"00",X"54",X"44",
		X"45",X"55",X"55",X"55",X"00",X"54",X"44",X"44",X"55",X"05",X"55",X"00",X"04",X"44",X"44",X"40",
		X"05",X"50",X"00",X"04",X"44",X"44",X"44",X"05",X"50",X"00",X"00",X"44",X"44",X"55",X"55",X"00",
		X"00",X"00",X"00",X"55",X"55",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F6",X"6F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"DC",X"F6",X"63",X"D6",X"66",X"66",X"66",
		X"6E",X"66",X"66",X"66",X"66",X"D3",X"66",X"00",X"D0",X"CC",X"CF",X"00",X"00",X"00",X"00",X"FF",
		X"0C",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"CC",X"FF",X"F0",X"00",X"0F",X"8F",
		X"FC",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"DC",X"6C",X"6F",X"FF",X"FF",X"88",
		X"89",X"6F",X"FF",X"0F",X"F0",X"00",X"00",X"00",X"00",X"DD",X"CF",X"FC",X"C8",X"88",X"8F",X"FC",
		X"6E",X"6F",X"66",X"F6",X"DF",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F8",X"8C",X"CC",X"CC",
		X"CC",X"CE",X"88",X"68",X"86",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"FF",X"CC",X"C6",
		X"6C",X"CC",X"98",X"69",X"86",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"CC",
		X"CC",X"CC",X"C9",X"69",X"98",X"6F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",
		X"CC",X"CC",X"CC",X"CC",X"C6",X"66",X"6F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"DF",X"CD",X"CC",X"CC",X"CC",X"C6",X"6B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",
		X"00",X"FD",X"FF",X"FC",X"CC",X"CC",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"CC",
		X"CC",X"6C",X"C6",X"6F",X"FF",X"FF",X"00",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F6",X"6F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"CC",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"DF",X"00",X"00",X"00",X"00",X"FF",
		X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"D0",X"DC",X"FF",X"F0",X"00",X"0F",X"6E",
		X"FC",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"0C",X"CC",X"6C",X"6F",X"FF",X"FF",X"CC",
		X"89",X"6F",X"FF",X"0F",X"F0",X"00",X"00",X"00",X"00",X"0C",X"CF",X"FC",X"CC",X"C6",X"6C",X"CC",
		X"88",X"6F",X"66",X"F6",X"DF",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FC",X"CC",X"CC",X"C8",
		X"88",X"CE",X"88",X"68",X"86",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"C8",X"88",
		X"8C",X"CC",X"98",X"69",X"86",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"CC",
		X"CC",X"CC",X"C9",X"69",X"98",X"6F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",
		X"CC",X"CC",X"CC",X"CC",X"C6",X"66",X"6F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"DF",X"CD",X"CC",X"CC",X"CC",X"C6",X"6B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",
		X"00",X"FD",X"FF",X"FC",X"CC",X"CC",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"CC",
		X"CC",X"6C",X"C6",X"6F",X"FF",X"FF",X"00",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F6",X"6F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"DD",X"F0",X"00",X"00",X"00",X"66",X"06",
		X"0C",X"60",X"60",X"66",X"00",X"00",X"00",X"00",X"00",X"CC",X"DF",X"00",X"00",X"00",X"00",X"FF",
		X"DC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"CC",X"FF",X"F0",X"00",X"0F",X"6E",
		X"FC",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"0C",X"CC",X"6C",X"6F",X"FF",X"FF",X"CC",
		X"69",X"8F",X"FF",X"0F",X"F0",X"00",X"00",X"00",X"0D",X"DC",X"CF",X"FC",X"CC",X"C6",X"6C",X"FC",
		X"6E",X"8F",X"88",X"F8",X"6F",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FC",X"CC",X"CC",X"CC",
		X"CC",X"CE",X"99",X"89",X"98",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"FF",X"CC",X"C6",
		X"6C",X"CC",X"99",X"89",X"98",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"CC",
		X"CC",X"CC",X"C9",X"69",X"99",X"6F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",
		X"CC",X"CC",X"CC",X"CC",X"C6",X"66",X"6F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"DF",X"CD",X"CC",X"CC",X"CC",X"C6",X"6B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",
		X"00",X"FD",X"FF",X"FC",X"CC",X"CC",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"CC",
		X"CC",X"6C",X"C6",X"6F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"44",
		X"04",X"D4",X"40",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"44",X"F4",X"F0",X"04",X"44",X"88",
		X"4C",X"00",X"04",X"44",X"40",X"40",X"00",X"00",X"00",X"44",X"00",X"04",X"44",X"4F",X"F4",X"44",
		X"00",X"C0",X"00",X"00",X"00",X"04",X"40",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"44",X"F4",
		X"4C",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"40",X"0C",X"C0",X"C0",X"00",X"C0",X"C0",
		X"CC",X"0E",X"44",X"44",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"04",X"CF",X"04",X"CE",
		X"44",X"BC",X"CC",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"CF",X"00",
		X"44",X"9C",X"CC",X"C0",X"C4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"CC",
		X"0C",X"CC",X"C0",X"4C",X"C4",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",
		X"CF",X"C4",X"CC",X"CC",X"04",X"44",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"FD",X"FC",X"FC",X"CC",X"C4",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"C0",
		X"CC",X"6C",X"00",X"0C",X"0C",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"50",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"05",X"00",X"00",X"00",X"00",X"50",
		X"00",X"05",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"50",X"05",X"00",X"55",X"05",X"00",
		X"05",X"00",X"00",X"50",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"55",
		X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"5F",X"55",X"0E",
		X"05",X"05",X"05",X"05",X"00",X"00",X"50",X"00",X"00",X"50",X"05",X"00",X"00",X"00",X"05",X"50",
		X"50",X"05",X"55",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"05",X"00",X"05",X"00",
		X"55",X"50",X"00",X"05",X"00",X"00",X"05",X"00",X"00",X"05",X"00",X"05",X"00",X"00",X"50",X"55",
		X"05",X"50",X"00",X"55",X"50",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"05",
		X"50",X"00",X"55",X"F0",X"05",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"50",
		X"05",X"05",X"05",X"05",X"50",X"5F",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"0E",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"00",X"EE",X"00",X"0E",
		X"00",X"00",X"00",X"E0",X"E0",X"00",X"00",X"00",X"0E",X"00",X"E0",X"00",X"E0",X"00",X"EE",X"00",
		X"0E",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"0E",X"0E",X"00",X"00",X"00",X"E0",X"EE",X"00",
		X"E0",X"00",X"E0",X"0E",X"00",X"00",X"E0",X"00",X"00",X"E0",X"0E",X"00",X"00",X"00",X"00",X"E0",
		X"E0",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"0E",X"00",
		X"0E",X"00",X"00",X"EE",X"00",X"0E",X"0E",X"00",X"E0",X"0E",X"00",X"0E",X"00",X"00",X"0E",X"00",
		X"0E",X"EE",X"0E",X"0E",X"E0",X"E0",X"00",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FB",X"BF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"DB",X"F6",X"63",X"D6",X"66",X"66",X"66",
		X"6E",X"66",X"66",X"66",X"66",X"D3",X"66",X"00",X"D0",X"BB",X"BF",X"00",X"00",X"00",X"00",X"FF",
		X"0B",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"BB",X"FF",X"F0",X"00",X"0F",X"BB",
		X"FB",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"DB",X"BB",X"BF",X"FF",X"FF",X"BB",
		X"BB",X"BF",X"FF",X"0F",X"F0",X"00",X"00",X"00",X"00",X"DD",X"BF",X"FB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BF",X"BB",X"FB",X"BF",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"22",X"B2",X"2B",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"FF",X"BB",X"BB",
		X"BB",X"BB",X"22",X"B2",X"2B",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"BB",
		X"BB",X"BB",X"B2",X"B2",X"22",X"BF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"BF",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",
		X"00",X"FB",X"FF",X"FB",X"BB",X"BB",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"BB",
		X"BB",X"BB",X"BB",X"BF",X"FF",X"FF",X"00",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F6",X"6F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"CC",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"DF",X"00",X"00",X"00",X"00",X"FF",
		X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"D0",X"DC",X"FF",X"F0",X"00",X"0F",X"6E",
		X"FC",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"0C",X"CC",X"6C",X"6F",X"FF",X"FF",X"C8",
		X"89",X"6F",X"FF",X"0F",X"F0",X"00",X"00",X"00",X"00",X"0C",X"CF",X"FC",X"CC",X"C6",X"6C",X"88",
		X"8C",X"6F",X"66",X"F6",X"DF",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FC",X"CC",X"C8",X"8C",
		X"CC",X"CE",X"88",X"68",X"86",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"86",
		X"6C",X"CC",X"98",X"69",X"86",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"8C",
		X"CC",X"CC",X"C9",X"69",X"98",X"6F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",
		X"CC",X"CC",X"CC",X"CC",X"C6",X"66",X"6F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"DF",X"CD",X"CC",X"CC",X"C8",X"86",X"6B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",
		X"00",X"FD",X"FF",X"FC",X"CC",X"CC",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"CC",
		X"CC",X"6C",X"C6",X"6F",X"FF",X"FF",X"00",X"00",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",
		X"54",X"20",X"28",X"43",X"29",X"20",X"31",X"39",X"38",X"34",X"2C",X"20",X"57",X"49",X"4C",X"4C",
		X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",
		X"20",X"49",X"4E",X"43",X"2E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"0F",X"00",X"40",X"00",X"00",X"00",X"40",X"0F",X"00",
		X"F0",X"04",X"40",X"00",X"00",X"00",X"44",X"00",X"F0",X"00",X"44",X"40",X"00",X"00",X"00",X"44",
		X"40",X"00",X"04",X"44",X"40",X"00",X"00",X"00",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"44",X"40",X"00",X"00",X"00",X"44",X"44",X"00",X"00",X"44",X"40",X"00",
		X"00",X"00",X"44",X"40",X"00",X"F0",X"04",X"40",X"00",X"00",X"00",X"44",X"00",X"F0",X"0F",X"00",
		X"40",X"00",X"00",X"00",X"40",X"0F",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"44",X"04",X"40",X"00",X"00",X"00",X"00",X"00",X"04",X"44",X"04",X"44",X"00",X"00",
		X"00",X"00",X"00",X"44",X"44",X"04",X"44",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"44",
		X"04",X"44",X"40",X"00",X"00",X"00",X"00",X"04",X"44",X"04",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"04",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"20",X"00",X"22",X"20",X"00",X"00",X"00",X"00",X"22",X"20",X"00",X"22",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"88",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"99",X"88",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"88",X"89",X"09",X"99",X"99",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"49",X"98",X"84",X"99",X"99",X"99",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"98",X"99",X"99",X"99",X"98",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"49",X"99",X"99",X"89",X"99",X"99",X"99",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"99",X"98",X"99",X"99",X"99",X"98",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"49",X"99",X"99",X"99",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"9A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"99",X"99",X"98",X"88",X"89",X"00",X"00",X"89",X"99",X"99",X"98",X"90",X"09",
		X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"99",X"99",X"99",X"88",X"88",
		X"9A",X"00",X"99",X"00",X"00",X"00",X"89",X"00",X"9A",X"00",X"00",X"00",X"00",X"00",X"66",X"DC",
		X"00",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"99",X"A9",X"90",X"00",X"00",X"08",X"9A",
		X"99",X"99",X"98",X"88",X"88",X"89",X"9C",X"C8",X"80",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"98",X"88",X"88",X"99",X"00",X"00",X"0A",X"89",X"99",X"99",X"99",X"99",X"99",X"99",X"CC",X"98",
		X"80",X"88",X"88",X"88",X"88",X"88",X"88",X"99",X"9A",X"98",X"88",X"88",X"88",X"88",X"89",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"89",X"98",X"D0",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"99",X"A9",X"99",X"CC",X"C9",X"99",X"99",X"98",X"88",X"99",X"99",X"99",X"98",X"88",X"88",X"9A",
		X"D0",X"49",X"99",X"99",X"99",X"98",X"88",X"88",X"88",X"9A",X"99",X"AA",X"A9",X"99",X"98",X"88",
		X"99",X"99",X"88",X"88",X"89",X"88",X"DA",X"A6",X"60",X"59",X"99",X"99",X"99",X"99",X"98",X"88",
		X"88",X"89",X"A9",X"99",X"99",X"99",X"88",X"99",X"99",X"88",X"88",X"88",X"88",X"98",X"DA",X"CC",
		X"C0",X"09",X"99",X"99",X"99",X"99",X"99",X"98",X"88",X"89",X"9A",X"99",X"99",X"99",X"99",X"99",
		X"98",X"88",X"88",X"88",X"88",X"89",X"C6",X"CC",X"00",X"00",X"00",X"00",X"0A",X"A9",X"99",X"99",
		X"88",X"88",X"9A",X"99",X"99",X"99",X"99",X"98",X"88",X"89",X"9A",X"A9",X"88",X"86",X"6C",X"00",
		X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"A9",X"99",X"98",X"88",X"9A",X"99",X"99",X"99",X"99",X"88",
		X"89",X"9A",X"AA",X"00",X"98",X"8C",X"C0",X"00",X"00",X"00",X"0A",X"A9",X"9D",X"99",X"AA",X"99",
		X"98",X"88",X"89",X"88",X"88",X"88",X"88",X"89",X"9A",X"A9",X"CD",X"99",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"99",X"CC",X"C8",X"9A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"09",X"CC",X"99",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"98",X"89",X"99",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A9",X"99",X"9A",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"99",X"99",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"88",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"99",X"88",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"88",X"89",X"09",X"99",X"99",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"49",X"98",X"84",X"99",X"99",X"99",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"98",X"99",X"99",X"99",X"98",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"49",X"99",X"99",X"89",X"99",X"99",X"99",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"99",X"98",X"99",X"99",X"99",X"98",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"49",X"99",X"99",X"99",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"9A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"99",X"99",X"98",X"88",X"89",X"00",X"00",X"89",X"99",X"99",X"98",X"90",X"09",
		X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"99",X"99",X"99",X"88",X"88",
		X"9A",X"00",X"99",X"00",X"00",X"00",X"89",X"00",X"9A",X"00",X"00",X"00",X"00",X"00",X"66",X"DC",
		X"00",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"99",X"A9",X"90",X"00",X"00",X"08",X"9A",
		X"99",X"99",X"98",X"88",X"88",X"89",X"9C",X"C8",X"80",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"98",X"88",X"88",X"99",X"00",X"00",X"0A",X"89",X"99",X"99",X"99",X"99",X"99",X"99",X"CC",X"98",
		X"80",X"88",X"88",X"88",X"88",X"88",X"88",X"99",X"9A",X"98",X"88",X"88",X"88",X"88",X"89",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"89",X"98",X"D0",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"99",X"A9",X"99",X"CC",X"C9",X"99",X"99",X"98",X"88",X"99",X"99",X"99",X"98",X"88",X"88",X"9A",
		X"D0",X"49",X"99",X"99",X"99",X"98",X"88",X"88",X"88",X"9A",X"99",X"AA",X"A9",X"99",X"98",X"88",
		X"99",X"99",X"88",X"88",X"89",X"88",X"DA",X"A6",X"60",X"59",X"99",X"99",X"99",X"99",X"98",X"88",
		X"88",X"89",X"A9",X"99",X"99",X"99",X"88",X"99",X"99",X"88",X"88",X"88",X"88",X"98",X"DA",X"CC",
		X"C0",X"09",X"99",X"99",X"99",X"99",X"99",X"98",X"88",X"89",X"9A",X"99",X"99",X"99",X"99",X"99",
		X"98",X"88",X"88",X"88",X"88",X"89",X"C6",X"CC",X"00",X"00",X"0A",X"AA",X"AA",X"A9",X"99",X"99",
		X"88",X"88",X"9A",X"99",X"99",X"99",X"99",X"98",X"88",X"89",X"AA",X"A9",X"88",X"86",X"6C",X"00",
		X"00",X"00",X"0A",X"A9",X"9D",X"99",X"A9",X"99",X"98",X"88",X"9A",X"99",X"99",X"99",X"99",X"88",
		X"89",X"A9",X"CD",X"99",X"A8",X"8C",X"C0",X"00",X"00",X"00",X"0A",X"99",X"CC",X"C8",X"9A",X"99",
		X"98",X"88",X"89",X"88",X"88",X"88",X"88",X"89",X"9A",X"A9",X"CC",X"99",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"98",X"89",X"99",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"A9",X"99",X"9A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"99",X"99",X"AA",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"AA",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"A8",X"89",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"98",X"89",X"94",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"89",X"99",X"99",X"09",X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"89",X"99",X"99",X"94",X"88",X"99",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"99",X"99",X"99",X"98",X"99",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"89",X"99",X"99",X"99",X"89",X"99",X"99",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"99",X"99",X"99",X"98",X"99",X"99",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"89",X"99",X"99",X"99",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A9",X"00",X"98",X"99",X"99",X"99",X"80",
		X"00",X"09",X"88",X"88",X"99",X"99",X"99",X"99",X"90",X"0C",X"D6",X"60",X"00",X"00",X"00",X"00",
		X"0A",X"90",X"09",X"80",X"00",X"00",X"09",X"90",X"0A",X"98",X"88",X"89",X"99",X"99",X"99",X"99",
		X"90",X"88",X"CC",X"99",X"88",X"88",X"88",X"99",X"99",X"9A",X"98",X"00",X"00",X"00",X"99",X"A9",
		X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"90",X"88",X"9C",X"C9",X"99",X"99",X"99",X"99",
		X"99",X"99",X"8A",X"00",X"00",X"09",X"98",X"88",X"88",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"90",X"D8",X"99",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"89",X"88",X"88",X"88",X"88",X"88",
		X"9A",X"99",X"98",X"88",X"88",X"88",X"88",X"88",X"80",X"DA",X"98",X"88",X"88",X"99",X"99",X"99",
		X"98",X"88",X"99",X"99",X"99",X"CC",X"C9",X"99",X"A9",X"98",X"88",X"88",X"88",X"88",X"88",X"88",
		X"80",X"66",X"AA",X"D8",X"89",X"88",X"88",X"89",X"99",X"98",X"88",X"99",X"99",X"AA",X"A9",X"9A",
		X"98",X"88",X"88",X"88",X"99",X"99",X"99",X"99",X"40",X"CC",X"CA",X"D8",X"98",X"88",X"88",X"88",
		X"89",X"99",X"98",X"89",X"99",X"99",X"99",X"A9",X"88",X"88",X"88",X"99",X"99",X"99",X"99",X"99",
		X"50",X"0C",X"C6",X"C9",X"88",X"88",X"88",X"88",X"88",X"99",X"99",X"99",X"99",X"99",X"9A",X"99",
		X"88",X"88",X"99",X"99",X"99",X"99",X"99",X"99",X"00",X"00",X"0C",X"66",X"88",X"89",X"AA",X"99",
		X"88",X"88",X"99",X"99",X"99",X"99",X"9A",X"98",X"88",X"89",X"99",X"99",X"AA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"CC",X"88",X"90",X"0A",X"AA",X"99",X"88",X"89",X"99",X"99",X"99",X"9A",X"98",
		X"88",X"99",X"99",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"A9",X"9D",X"C9",
		X"AA",X"99",X"88",X"88",X"88",X"88",X"89",X"88",X"88",X"99",X"9A",X"A9",X"9D",X"99",X"AA",X"00",
		X"00",X"00",X"00",X"00",X"00",X"A9",X"9C",X"C9",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"AA",X"98",X"CC",X"C9",X"9A",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"99",X"99",
		X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A9",X"99",X"88",X"99",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"A9",X"99",X"9A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"A8",X"89",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"98",X"89",X"94",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"89",X"99",X"99",X"09",X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"89",X"99",X"99",X"94",X"88",X"99",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"99",X"99",X"99",X"98",X"99",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"89",X"99",X"99",X"99",X"89",X"99",X"99",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"99",X"99",X"99",X"98",X"99",X"99",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"89",X"99",X"99",X"99",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A9",X"00",X"98",X"99",X"99",X"99",X"80",
		X"00",X"09",X"88",X"88",X"99",X"99",X"99",X"99",X"90",X"0C",X"D6",X"60",X"00",X"00",X"00",X"00",
		X"0A",X"90",X"09",X"80",X"00",X"00",X"09",X"90",X"0A",X"98",X"88",X"89",X"99",X"99",X"99",X"99",
		X"90",X"88",X"CC",X"99",X"88",X"88",X"88",X"99",X"99",X"9A",X"98",X"00",X"00",X"00",X"99",X"A9",
		X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"90",X"88",X"9C",X"C9",X"99",X"99",X"99",X"99",
		X"99",X"99",X"8A",X"00",X"00",X"09",X"98",X"88",X"88",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"90",X"D8",X"99",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"89",X"88",X"88",X"88",X"88",X"88",
		X"9A",X"99",X"98",X"88",X"88",X"88",X"88",X"88",X"80",X"DA",X"98",X"88",X"88",X"99",X"99",X"99",
		X"98",X"88",X"99",X"99",X"99",X"CC",X"C9",X"99",X"A9",X"98",X"88",X"88",X"88",X"88",X"88",X"88",
		X"80",X"66",X"AA",X"D8",X"89",X"88",X"88",X"89",X"99",X"98",X"88",X"99",X"99",X"AA",X"A9",X"9A",
		X"98",X"88",X"88",X"88",X"99",X"99",X"99",X"99",X"40",X"CC",X"CA",X"D8",X"98",X"88",X"88",X"88",
		X"89",X"99",X"98",X"89",X"99",X"99",X"99",X"A9",X"88",X"88",X"88",X"99",X"99",X"99",X"99",X"99",
		X"50",X"0C",X"C6",X"C9",X"88",X"88",X"88",X"88",X"88",X"99",X"99",X"99",X"99",X"99",X"9A",X"99",
		X"88",X"88",X"99",X"99",X"99",X"99",X"99",X"99",X"00",X"00",X"0C",X"66",X"88",X"89",X"AA",X"A9",
		X"88",X"88",X"99",X"99",X"99",X"99",X"9A",X"98",X"88",X"89",X"99",X"99",X"AA",X"AA",X"AA",X"00",
		X"00",X"00",X"00",X"CC",X"88",X"A9",X"9D",X"C9",X"A9",X"88",X"89",X"99",X"99",X"99",X"9A",X"98",
		X"88",X"99",X"99",X"A9",X"9D",X"99",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"A9",X"9C",X"C9",
		X"AA",X"99",X"88",X"88",X"88",X"88",X"89",X"88",X"88",X"99",X"9A",X"98",X"CC",X"C9",X"9A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"99",X"99",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A9",X"99",X"88",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"A9",X"99",X"9A",X"00",X"00",
		X"00",X"0F",X"F0",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"F0",X"00",X"FF",X"44",X"44",X"0F",X"00",
		X"0F",X"44",X"44",X"40",X"00",X"00",X"42",X"44",X"40",X"00",X"00",X"44",X"24",X"40",X"00",X"00",
		X"04",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"F0",X"00",X"0F",X"FF",X"FF",
		X"00",X"00",X"F4",X"00",X"F0",X"00",X"44",X"40",X"F0",X"04",X"24",X"44",X"F0",X"04",X"24",X"44",
		X"F0",X"04",X"44",X"44",X"00",X"00",X"40",X"40",X"00",X"0F",X"FF",X"00",X"00",X"FF",X"F0",X"F0",
		X"00",X"FF",X"44",X"4F",X"00",X"04",X"44",X"44",X"00",X"04",X"24",X"44",X"00",X"00",X"42",X"40",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"F0",X"00",X"00",X"FF",X"0F",X"00",X"00",X"44",X"0F",
		X"00",X"04",X"24",X"4F",X"00",X"04",X"24",X"40",X"00",X"04",X"44",X"40",X"00",X"00",X"44",X"00",
		X"00",X"0F",X"F0",X"00",X"FF",X"44",X"00",X"04",X"44",X"40",X"04",X"24",X"40",X"00",X"44",X"00",
		X"0F",X"FF",X"00",X"04",X"40",X"F0",X"42",X"44",X"40",X"42",X"44",X"40",X"44",X"44",X"40",X"04",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"44",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"44",X"44",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4E",
		X"44",X"4E",X"40",X"00",X"00",X"00",X"00",X"00",X"04",X"4E",X"45",X"4E",X"44",X"00",X"00",X"00",
		X"00",X"00",X"00",X"4E",X"45",X"4E",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"45",X"4E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"4E",X"4E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",
		X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"EE",X"EE",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0D",X"CE",X"44",X"4E",X"40",X"00",X"00",X"00",X"00",X"00",X"0D",X"CE",X"45",X"4E",
		X"44",X"00",X"00",X"00",X"00",X"00",X"0C",X"CE",X"45",X"4E",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"45",X"4E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"4E",X"4E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"44",X"44",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"0E",X"EE",X"EE",
		X"00",X"00",X"00",X"00",X"D6",X"DD",X"DD",X"CE",X"44",X"4E",X"40",X"00",X"00",X"00",X"6D",X"DD",
		X"DD",X"CE",X"45",X"4E",X"44",X"00",X"00",X"00",X"D9",X"CC",X"CC",X"CE",X"45",X"4E",X"40",X"00",
		X"00",X"00",X"0D",X"00",X"00",X"0E",X"45",X"4E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",
		X"4E",X"4E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"44",X"44",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"44",X"44",X"00",X"00",X"0D",X"D0",X"00",X"00",
		X"00",X"0E",X"EE",X"EE",X"00",X"00",X"DD",X"6D",X"DD",X"DD",X"DD",X"CE",X"44",X"4E",X"40",X"00",
		X"6D",X"DD",X"DD",X"DD",X"DD",X"CE",X"45",X"4E",X"44",X"00",X"DD",X"6C",X"CC",X"CC",X"CC",X"CE",
		X"45",X"4E",X"40",X"00",X"0D",X"D0",X"00",X"00",X"00",X"0E",X"45",X"4E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"4E",X"4E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"44",X"44",
		X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"05",X"E5",X"00",X"00",X"00",X"4E",X"4E",
		X"40",X"00",X"00",X"0E",X"4E",X"00",X"00",X"00",X"0E",X"EE",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"05",X"E5",X"00",X"00",X"00",X"6E",X"4E",X"40",X"00",X"00",X"0E",X"4E",X"00",X"00",
		X"00",X"0E",X"EE",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"05",X"E5",X"00",X"00",X"DD",
		X"6E",X"4E",X"40",X"00",X"00",X"0E",X"4E",X"00",X"00",X"00",X"0E",X"EE",X"00",X"00",X"00",X"00",
		X"40",X"00",X"60",X"00",X"05",X"E5",X"00",X"DD",X"DD",X"6E",X"4E",X"40",X"60",X"00",X"0E",X"4E",
		X"00",X"00",X"00",X"0E",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"9E",X"5E",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"44",X"50",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"55",X"54",X"5E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"55",X"45",X"50",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"0E",X"5E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"E5",X"75",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"5E",X"55",X"55",
		X"50",X"00",X"00",X"00",X"00",X"00",X"05",X"50",X"EE",X"EE",X"E0",X"54",X"00",X"00",X"00",X"00",
		X"00",X"55",X"00",X"E5",X"E5",X"E0",X"05",X"50",X"00",X"00",X"00",X"05",X"55",X"00",X"E5",X"55",
		X"E0",X"05",X"55",X"00",X"00",X"00",X"E4",X"5E",X"00",X"5E",X"54",X"50",X"0E",X"54",X"E0",X"00",
		X"00",X"45",X"E5",X"00",X"5E",X"55",X"40",X"05",X"E5",X"40",X"00",X"05",X"54",X"EE",X"00",X"EE",
		X"54",X"E0",X"0E",X"E4",X"55",X"00",X"E4",X"E5",X"50",X"00",X"0E",X"EE",X"00",X"00",X"55",X"E4",
		X"E0",X"55",X"EE",X"50",X"00",X"0E",X"4E",X"00",X"00",X"5E",X"E5",X"50",X"45",X"E0",X"50",X"00",
		X"05",X"55",X"00",X"00",X"50",X"E5",X"40",X"55",X"E0",X"E0",X"00",X"55",X"E4",X"50",X"00",X"E0",
		X"E5",X"50",X"04",X"50",X"E0",X"0E",X"5E",X"E0",X"5E",X"00",X"E0",X"54",X"00",X"0E",X"50",X"00",
		X"05",X"EE",X"4E",X"05",X"00",X"00",X"50",X"00",X"00",X"50",X"00",X"00",X"50",X"4E",X"50",X"00",
		X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"40",X"E0",X"40",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"B4",X"E4",X"B0",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"0B",X"5B",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E5",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"55",
		X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"5E",X"55",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E5",X"50",X"0F",X"4F",X"EE",X"B0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E5",X"E0",X"0E",X"E5",X"E5",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"5E",
		X"00",X"0E",X"55",X"4E",X"E5",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"E5",X"00",X"0A",X"AE",
		X"55",X"05",X"50",X"00",X"00",X"00",X"00",X"04",X"E5",X"00",X"00",X"EA",X"4A",X"5E",X"0E",X"5E",
		X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"45",X"54",X"A0",X"00",X"55",X"00",X"00",X"00",
		X"00",X"05",X"00",X"00",X"0E",X"EE",X"A5",X"E0",X"00",X"54",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"EB",X"EE",X"40",X"05",X"E5",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B5",
		X"BE",X"E0",X"00",X"05",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"55",X"BE",X"00",X"00",
		X"40",X"E4",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"05",X"4B",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"5B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"40",X"50",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"EE",X"5E",X"00",
		X"55",X"45",X"50",X"0E",X"55",X"80",X"00",X"00",X"00",X"0E",X"EE",X"EE",X"EE",X"05",X"E5",X"00",
		X"E5",X"54",X"90",X"00",X"00",X"00",X"E0",X"0E",X"00",X"00",X"0E",X"EE",X"55",X"0E",X"55",X"5B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B4",X"AE",X"E5",X"54",X"55",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E4",X"5E",X"54",X"E5",X"50",X"4E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B4",X"EE",X"EB",X"55",X"50",X"E5",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"45",X"E4",X"BE",
		X"5E",X"00",X"05",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"E0",X"00",X"00",X"0E",
		X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E5",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"54",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"E5",X"50",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"05",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E5",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",
		X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"50",X"05",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"55",X"4E",X"50",X"0E",X"55",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"E5",X"00",X"05",X"54",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"EE",X"55",
		X"EE",X"55",X"5B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"AE",X"E5",X"54",X"55",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"5B",X"5E",X"5B",X"E5",X"50",X"4E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"BB",X"EE",X"EB",X"55",X"50",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"4B",X"EB",X"BE",X"5E",X"00",X"05",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"E0",
		X"00",X"00",X"0E",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"05",
		X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"0E",X"55",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"E5",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"05",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"5E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"50",X"00",X"00",X"00",
		X"40",X"00",X"E5",X"00",X"00",X"00",X"E4",X"50",X"05",X"00",X"00",X"00",X"04",X"00",X"05",X"00",
		X"00",X"04",X"BE",X"55",X"EE",X"00",X"00",X"BB",X"EB",X"E5",X"50",X"00",X"00",X"0E",X"BE",X"E5",
		X"5E",X"59",X"00",X"0B",X"40",X"E5",X"EE",X"5E",X"00",X"00",X"00",X"00",X"5E",X"5B",X"00",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"0E",X"E5",X"00",
		X"00",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"00",X"05",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"50",X"00",X"00",X"00",X"00",X"00",X"EE",X"50",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"00",X"04",X"BE",X"EE",X"00",X"00",X"00",X"BB",X"EB",X"E5",X"50",X"00",X"00",X"0E",X"BE",X"E5",
		X"5E",X"59",X"00",X"0B",X"50",X"EE",X"EE",X"5E",X"00",X"00",X"00",X"00",X"5E",X"5B",X"00",X"00",
		X"00",X"E5",X"E0",X"00",X"00",X"00",X"0E",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"E0",X"05",X"BE",X"00",
		X"00",X"00",X"E0",X"00",X"EE",X"50",X"00",X"EE",X"00",X"00",X"0E",X"55",X"0E",X"E0",X"00",X"00",
		X"00",X"E5",X"50",X"00",X"00",X"00",X"00",X"E5",X"E9",X"00",X"00",X"00",X"00",X"E0",X"5B",X"90",
		X"00",X"00",X"EE",X"00",X"09",X"E0",X"00",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0B",X"00",X"0E",X"00",X"00",X"00",X"05",X"BE",X"00",X"E0",X"00",X"00",X"00",
		X"EE",X"50",X"E0",X"00",X"00",X"00",X"0E",X"55",X"E0",X"00",X"00",X"0E",X"00",X"E5",X"50",X"00",
		X"00",X"00",X"EE",X"E5",X"E9",X"00",X"00",X"00",X"00",X"00",X"5B",X"90",X"00",X"00",X"00",X"00",
		X"09",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"F0",X"00",X"00",X"0F",X"FC",X"CF",X"00",X"00",X"FC",X"CC",X"CF",X"00",X"00",X"FC",X"CD",X"CC",
		X"F0",X"00",X"0F",X"CC",X"CF",X"00",X"00",X"00",X"FC",X"F0",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"F0",X"00",X"00",X"FF",X"CD",X"CF",X"00",X"00",
		X"CC",X"FC",X"FF",X"F0",X"00",X"CD",X"F0",X"0C",X"DF",X"00",X"FC",X"FD",X"0C",X"CC",X"00",X"0F",
		X"F0",X"0F",X"F0",X"00",X"FC",X"CF",X"CC",X"CF",X"00",X"FC",X"CD",X"FC",X"CF",X"00",X"0F",X"CF",
		X"FC",X"F0",X"00",X"00",X"FD",X"F0",X"00",X"00",X"FF",X"CF",X"CF",X"00",X"00",X"CF",X"F0",X"F0",
		X"0F",X"00",X"DF",X"00",X"00",X"FD",X"00",X"CF",X"0D",X"0F",X"CC",X"00",X"FF",X"00",X"00",X"FF",
		X"00",X"FC",X"F0",X"0F",X"CF",X"00",X"FC",X"FF",X"0F",X"CF",X"00",X"0F",X"CD",X"FC",X"F0",X"00",
		X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",
		X"00",X"00",X"05",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"0E",
		X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0D",X"D0",X"00",X"D0",X"0D",X"00",
		X"D0",X"0D",X"00",X"D0",X"0D",X"00",X"D0",X"0D",X"00",X"D0",X"0D",X"00",X"0D",X"D0",X"00",X"0D",
		X"00",X"00",X"DD",X"00",X"00",X"0D",X"00",X"00",X"0D",X"00",X"00",X"0D",X"00",X"00",X"0D",X"00",
		X"00",X"DD",X"D0",X"00",X"0D",X"D0",X"00",X"D0",X"0D",X"00",X"00",X"0D",X"00",X"00",X"D0",X"00",
		X"0D",X"00",X"00",X"D0",X"00",X"00",X"DD",X"DD",X"00",X"0D",X"D0",X"00",X"D0",X"0D",X"00",X"00",
		X"0D",X"00",X"0D",X"D0",X"00",X"00",X"0D",X"00",X"D0",X"0D",X"00",X"0D",X"D0",X"00",X"00",X"D0",
		X"00",X"D0",X"D0",X"00",X"D0",X"D0",X"00",X"DD",X"DD",X"00",X"00",X"D0",X"00",X"00",X"D0",X"00",
		X"00",X"D0",X"00",X"DD",X"D0",X"00",X"D0",X"00",X"00",X"DD",X"D0",X"00",X"00",X"0D",X"00",X"00",
		X"0D",X"00",X"D0",X"0D",X"00",X"0D",X"D0",X"00",X"0D",X"D0",X"00",X"D0",X"00",X"00",X"D0",X"00",
		X"00",X"DD",X"D0",X"00",X"D0",X"0D",X"00",X"D0",X"0D",X"00",X"0D",X"D0",X"00",X"DD",X"DD",X"00",
		X"00",X"0D",X"00",X"00",X"0D",X"00",X"00",X"D0",X"00",X"0D",X"00",X"00",X"0D",X"00",X"00",X"0D",
		X"00",X"00",X"0D",X"D0",X"00",X"D0",X"0D",X"00",X"0D",X"D0",X"00",X"D0",X"0D",X"00",X"D0",X"0D",
		X"00",X"D0",X"0D",X"00",X"0D",X"D0",X"00",X"0D",X"D0",X"00",X"D0",X"0D",X"00",X"D0",X"0D",X"00",
		X"0D",X"DD",X"00",X"00",X"0D",X"00",X"D0",X"0D",X"00",X"0D",X"D0",X"00",X"00",X"DD",X"00",X"0D",
		X"CC",X"C0",X"0C",X"CC",X"00",X"00",X"C0",X"00",X"00",X"0F",X"F0",X"0D",X"C0",X"00",X"DC",X"CC",
		X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"80",X"00",X"00",X"86",X"66",X"66",X"68",
		X"00",X"08",X"89",X"99",X"90",X"00",X"06",X"66",X"88",X"80",X"00",X"66",X"66",X"A6",X"88",X"00",
		X"06",X"86",X"A6",X"80",X"00",X"06",X"86",X"96",X"80",X"00",X"06",X"86",X"96",X"80",X"00",X"06",
		X"96",X"A6",X"80",X"00",X"06",X"96",X"A6",X"80",X"00",X"06",X"A6",X"96",X"80",X"00",X"06",X"86",
		X"86",X"80",X"00",X"00",X"00",X"B0",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"50",X"00",X"00",X"60",
		X"00",X"5B",X"00",X"06",X"0B",X"00",X"00",X"00",X"60",X"00",X"05",X"00",X"00",X"60",X"00",X"00",
		X"00",X"66",X"60",X"0B",X"50",X"E0",X"56",X"00",X"00",X"00",X"06",X"88",X"00",X"BE",X"0B",X"00",
		X"0B",X"00",X"00",X"00",X"00",X"0E",X"22",X"B5",X"50",X"00",X"00",X"00",X"00",X"00",X"05",X"42",
		X"50",X"00",X"06",X"60",X"06",X"00",X"05",X"B2",X"BD",X"5B",X"00",X"66",X"80",X"66",X"60",X"50",
		X"5B",X"DB",X"B0",X"66",X"66",X"A0",X"06",X"66",X"60",X"05",X"52",X"50",X"00",X"68",X"00",X"06",
		X"80",X"00",X"E0",X"D2",X"2B",X"00",X"0A",X"00",X"08",X"00",X"00",X"0B",X"45",X"05",X"B0",X"00",
		X"00",X"00",X"00",X"60",X"5B",X"0E",X"00",X"50",X"00",X"00",X"00",X"06",X"60",X"50",X"00",X"00",
		X"00",X"60",X"00",X"09",X"00",X"0B",X"50",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"06",
		X"68",X"00",X"00",X"0B",X"00",X"00",X"00",X"06",X"66",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"0B",X"00",X"00",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"0B",
		X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"6A",X"00",X"86",X"66",X"80",X"08",X"99",X"00",X"66",X"88",
		X"80",X"A6",X"68",X"00",X"06",X"68",X"00",X"06",X"68",X"00",X"06",X"68",X"00",X"00",X"00",X"00",
		X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"60",X"00",X"00",X"06",X"00",X"06",
		X"80",X"00",X"0B",X"00",X"60",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"02",X"40",X"00",
		X"00",X"66",X"04",X"B2",X"00",X"06",X"80",X"08",X"60",X"0B",X"B0",X"50",X"00",X"00",X"00",X"50",
		X"40",X"00",X"00",X"06",X"05",X"00",X"04",X"00",X"60",X"00",X"00",X"0A",X"60",X"00",X"00",X"00",
		X"00",X"66",X"60",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"50",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"28",X"43",X"29",X"20",X"31",X"39",
		X"38",X"34",X"2C",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",
		X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"00",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9E",X"5E",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"54",X"45",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"54",X"55",X"5E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"55",X"45",X"50",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"5E",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"E5",X"75",X"EE",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"55",X"55",X"5E",X"55",X"50",X"00",X"00",X"00",X"00",X"00",X"04",X"50",X"EE",
		X"EE",X"E0",X"55",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"E5",X"E5",X"E0",X"05",X"50",X"00",
		X"00",X"00",X"05",X"55",X"00",X"E5",X"55",X"E0",X"05",X"55",X"00",X"00",X"00",X"E4",X"5E",X"00",
		X"54",X"5E",X"50",X"0E",X"54",X"E0",X"00",X"00",X"45",X"E5",X"00",X"45",X"5E",X"50",X"05",X"E5",
		X"40",X"00",X"05",X"54",X"EE",X"00",X"E4",X"5E",X"E0",X"0E",X"E4",X"55",X"00",X"E4",X"E5",X"50",
		X"00",X"0E",X"EE",X"00",X"00",X"55",X"E4",X"E0",X"55",X"EE",X"50",X"00",X"0E",X"4E",X"00",X"00",
		X"5E",X"E5",X"50",X"45",X"E0",X"50",X"00",X"05",X"55",X"00",X"00",X"50",X"E5",X"40",X"55",X"E0",
		X"E0",X"00",X"54",X"E5",X"50",X"00",X"E0",X"E5",X"50",X"04",X"50",X"E0",X"0E",X"50",X"EE",X"5E",
		X"00",X"E0",X"54",X"00",X"00",X"50",X"00",X"05",X"0E",X"4E",X"E5",X"00",X"00",X"5E",X"00",X"00",
		X"50",X"00",X"00",X"5E",X"40",X"50",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"40",X"E0",
		X"40",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"B4",X"E4",X"B0",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"0B",X"5B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"05",X"5E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"54",X"55",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",
		X"E5",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"EE",X"F4",X"F0",X"05",
		X"5E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"5E",X"5E",X"E0",X"0E",X"5E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"5E",X"E4",X"55",X"E0",X"00",X"E5",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"05",X"50",X"55",X"EA",X"A0",X"00",X"5E",X"40",X"00",X"00",X"00",X"00",X"00",X"E5",
		X"E0",X"E5",X"A4",X"AE",X"00",X"00",X"5E",X"40",X"00",X"00",X"00",X"00",X"55",X"00",X"0A",X"45",
		X"54",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"45",X"00",X"0E",X"5A",X"EE",X"E0",X"00",
		X"00",X"50",X"00",X"00",X"00",X"0E",X"5E",X"50",X"04",X"EE",X"BE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"50",X"00",X"0E",X"EB",X"5B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4E",
		X"04",X"00",X"00",X"EB",X"55",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B4",X"50",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B5",X"0B",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"05",X"04",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"55",X"E0",X"05",X"54",X"55",X"00",X"E5",X"EE",X"00",X"00",
		X"00",X"00",X"09",X"45",X"5E",X"00",X"5E",X"50",X"EE",X"EE",X"EE",X"E0",X"00",X"00",X"00",X"B5",
		X"55",X"E0",X"55",X"EE",X"E0",X"00",X"00",X"E0",X"0E",X"00",X"00",X"00",X"0E",X"55",X"45",X"5E",
		X"EA",X"4B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E4",X"05",X"5E",X"45",X"E5",X"4E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5E",X"05",X"55",X"BE",X"EE",X"4B",X"00",X"00",X"00",
		X"00",X"00",X"00",X"05",X"50",X"00",X"E5",X"EB",X"4E",X"54",X"00",X"00",X"00",X"00",X"00",X"00",
		X"45",X"E0",X"00",X"00",X"0E",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"5E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"45",X"50",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"05",X"5E",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",
		X"5E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"50",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"50",X"05",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"55",X"E0",X"05",X"E4",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"45",X"50",X"00",X"5E",X"50",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"B5",X"55",X"EE",X"55",X"EE",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"55",X"45",X"5E",X"EA",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E4",
		X"05",X"5E",X"B5",X"E5",X"B5",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"05",X"55",X"BE",
		X"EE",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"50",X"00",X"E5",X"EB",X"BE",X"B4",X"00",
		X"00",X"00",X"00",X"00",X"00",X"05",X"E0",X"00",X"00",X"0E",X"BB",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"05",X"50",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",
		X"55",X"E0",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5E",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"50",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"50",X"05",X"00",X"00",X"00",X"05",X"E0",X"00",X"40",X"00",X"00",X"05",X"00",X"54",
		X"E0",X"00",X"00",X"05",X"00",X"04",X"00",X"00",X"00",X"0E",X"E5",X"5E",X"B4",X"00",X"00",X"00",
		X"55",X"EB",X"EB",X"B0",X"09",X"5E",X"55",X"EE",X"BE",X"00",X"0E",X"5E",X"E5",X"E0",X"4B",X"00",
		X"0B",X"5E",X"50",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"00",X"05",X"EE",X"00",X"00",X"00",X"00",X"0E",X"50",X"00",X"00",X"00",X"00",X"00",
		X"E5",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"5E",
		X"E0",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"0E",X"EE",X"B4",X"00",X"00",X"00",
		X"55",X"EB",X"EB",X"B0",X"09",X"5E",X"55",X"EE",X"BE",X"00",X"0E",X"5E",X"EE",X"E0",X"5B",X"00",
		X"0B",X"5E",X"50",X"00",X"00",X"00",X"00",X"00",X"E5",X"E0",X"00",X"00",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"0B",X"00",X"E0",X"00",X"00",X"0E",X"B5",X"00",X"0E",X"E0",X"00",X"5E",X"E0",X"00",
		X"00",X"EE",X"05",X"5E",X"00",X"00",X"00",X"00",X"55",X"E0",X"00",X"00",X"00",X"09",X"E5",X"E0",
		X"00",X"00",X"00",X"9B",X"50",X"E0",X"00",X"00",X"00",X"E9",X"00",X"0E",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"0B",X"00",
		X"00",X"00",X"E0",X"0E",X"B5",X"00",X"00",X"00",X"E0",X"5E",X"E0",X"00",X"00",X"00",X"E5",X"5E",
		X"00",X"00",X"00",X"00",X"55",X"E0",X"0E",X"00",X"00",X"09",X"E5",X"EE",X"E0",X"00",X"00",X"9B",
		X"50",X"00",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"44",X"00",X"00",X"00",X"00",X"05",X"55",X"45",X"55",X"00",X"00",X"00",X"55",
		X"E5",X"54",X"55",X"50",X"00",X"00",X"55",X"E5",X"45",X"E5",X"50",X"00",X"00",X"E5",X"EE",X"EE",
		X"E5",X"E0",X"00",X"00",X"0E",X"5E",X"EE",X"5E",X"00",X"00",X"00",X"00",X"EE",X"EE",X"E0",X"00",
		X"00",X"00",X"0D",X"CD",X"DD",X"CD",X"00",X"00",X"00",X"06",X"66",X"66",X"66",X"00",X"00",X"00",
		X"C6",X"66",X"66",X"66",X"C0",X"00",X"00",X"66",X"66",X"C6",X"66",X"60",X"00",X"00",X"66",X"C4",
		X"44",X"C6",X"60",X"00",X"00",X"CC",X"9C",X"6C",X"9C",X"C0",X"00",X"00",X"09",X"C6",X"66",X"C9",
		X"00",X"00",X"00",X"0E",X"C6",X"66",X"CE",X"00",X"00",X"00",X"00",X"C6",X"66",X"C0",X"00",X"00",
		X"00",X"00",X"66",X"66",X"60",X"00",X"00",X"00",X"00",X"66",X"66",X"60",X"00",X"00",X"00",X"00",
		X"66",X"66",X"60",X"00",X"00",X"00",X"00",X"09",X"09",X"00",X"00",X"00",X"00",X"00",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"00",X"00",
		X"00",X"00",X"00",X"55",X"E5",X"50",X"00",X"00",X"00",X"00",X"5E",X"4E",X"50",X"00",X"00",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"07",X"54",X"55",X"00",X"00",X"07",X"77",X"07",
		X"75",X"44",X"50",X"00",X"00",X"77",X"77",X"75",X"45",X"50",X"00",X"00",X"47",X"75",X"55",X"50",
		X"00",X"00",X"00",X"07",X"75",X"55",X"40",X"00",X"00",X"00",X"00",X"77",X"55",X"50",X"00",X"00",
		X"00",X"00",X"0D",X"DD",X"D0",X"00",X"00",X"00",X"00",X"DD",X"66",X"68",X"00",X"00",X"00",X"06",
		X"66",X"68",X"66",X"80",X"00",X"00",X"66",X"66",X"C0",X"06",X"60",X"00",X"00",X"C6",X"6C",X"40",
		X"00",X"66",X"00",X"00",X"00",X"94",X"46",X"C0",X"66",X"00",X"00",X"0C",X"0C",X"66",X"60",X"77",
		X"00",X"00",X"07",X"00",X"66",X"85",X"77",X"50",X"00",X"70",X"00",X"66",X"85",X"99",X"40",X"00",
		X"00",X"00",X"66",X"84",X"55",X"40",X"00",X"00",X"00",X"6C",X"84",X"44",X"40",X"00",X"00",X"06",
		X"6C",X"84",X"44",X"40",X"00",X"00",X"00",X"C5",X"09",X"00",X"00",X"00",X"00",X"00",X"77",X"07",
		X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"70",X"00",X"00",X"00",X"07",X"00",X"00",X"04",X"50",
		X"00",X"00",X"74",X"00",X"00",X"05",X"00",X"00",X"44",X"04",X"00",X"00",X"55",X"00",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"07",X"54",X"55",X"00",X"00",X"07",X"77",X"07",X"75",
		X"44",X"50",X"00",X"00",X"77",X"77",X"75",X"45",X"50",X"00",X"00",X"47",X"75",X"55",X"50",X"00",
		X"00",X"00",X"07",X"75",X"55",X"40",X"00",X"00",X"00",X"00",X"77",X"55",X"50",X"00",X"00",X"00",
		X"00",X"0D",X"DD",X"D0",X"00",X"00",X"00",X"00",X"DD",X"66",X"C0",X"00",X"00",X"00",X"06",X"66",
		X"86",X"68",X"00",X"00",X"00",X"66",X"66",X"C0",X"C6",X"80",X"00",X"00",X"C6",X"6C",X"40",X"0C",
		X"60",X"00",X"00",X"00",X"04",X"46",X"06",X"C0",X"00",X"00",X"00",X"0C",X"66",X"66",X"00",X"00",
		X"00",X"00",X"00",X"67",X"70",X"00",X"00",X"00",X"00",X"00",X"57",X"70",X"00",X"00",X"00",X"00",
		X"00",X"58",X"85",X"00",X"00",X"00",X"00",X"00",X"45",X"54",X"00",X"00",X"00",X"00",X"00",X"44",
		X"44",X"00",X"00",X"00",X"00",X"00",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",
		X"00",X"00",X"07",X"40",X"00",X"00",X"00",X"00",X"04",X"40",X"40",X"00",X"00",X"00",X"00",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"75",X"45",X"50",X"00",X"00",X"77",X"70",X"77",X"54",X"45",
		X"00",X"00",X"07",X"77",X"77",X"54",X"55",X"00",X"00",X"04",X"77",X"55",X"55",X"00",X"00",X"00",
		X"00",X"77",X"55",X"54",X"00",X"00",X"00",X"00",X"07",X"75",X"55",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"DD",X"00",X"00",X"00",X"00",X"0D",X"D6",X"60",X"00",X"00",X"00",X"00",X"66",X"6C",X"60",
		X"00",X"00",X"00",X"06",X"66",X"CC",X"60",X"00",X"00",X"00",X"0C",X"66",X"C6",X"60",X"00",X"00",
		X"00",X"00",X"00",X"66",X"C0",X"00",X"00",X"00",X"00",X"06",X"6C",X"86",X"00",X"00",X"00",X"00",
		X"66",X"08",X"C6",X"00",X"00",X"00",X"07",X"70",X"0C",X"66",X"00",X"00",X"00",X"57",X"70",X"06",
		X"66",X"00",X"00",X"00",X"59",X"95",X"0C",X"66",X"60",X"00",X"00",X"45",X"54",X"09",X"00",X"77",
		X"00",X"00",X"44",X"44",X"57",X"00",X"07",X"00",X"00",X"44",X"44",X"00",X"00",X"0E",X"74",X"40",
		X"00",X"00",X"50",X"00",X"00",X"74",X"00",X"00",X"74",X"00",X"00",X"00",X"04",X"50",X"04",X"04",
		X"00",X"00",X"00",X"00",X"40",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"40",
		X"00",X"00",X"00",X"00",X"05",X"77",X"77",X"50",X"00",X"00",X"00",X"54",X"00",X"70",X"55",X"00",
		X"00",X"00",X"47",X"77",X"77",X"74",X"00",X"00",X"00",X"05",X"77",X"57",X"50",X"00",X"00",X"00",
		X"00",X"57",X"75",X"00",X"00",X"00",X"00",X"0D",X"D7",X"7D",X"D0",X"00",X"00",X"00",X"C6",X"CD",
		X"DC",X"6C",X"00",X"00",X"00",X"66",X"66",X"66",X"66",X"00",X"00",X"00",X"C7",X"75",X"57",X"7C",
		X"00",X"00",X"00",X"07",X"48",X"84",X"70",X"00",X"00",X"00",X"00",X"45",X"54",X"00",X"00",X"00",
		X"00",X"00",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"00",
		X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"70",
		X"00",X"00",X"00",X"00",X"00",X"07",X"70",X"00",X"00",X"00",X"00",X"00",X"07",X"70",X"00",X"00",
		X"00",X"00",X"00",X"57",X"75",X"00",X"00",X"00",X"00",X"00",X"44",X"54",X"00",X"00",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"75",X"45",X"50",X"00",X"00",X"07",X"70",X"77",
		X"54",X"55",X"00",X"00",X"00",X"77",X"77",X"55",X"55",X"00",X"00",X"00",X"47",X"75",X"54",X"00",
		X"00",X"00",X"00",X"00",X"77",X"55",X"00",X"00",X"00",X"00",X"00",X"0D",X"DD",X"00",X"00",X"00",
		X"00",X"00",X"D6",X"66",X"60",X"00",X"00",X"00",X"96",X"66",X"80",X"C6",X"00",X"00",X"00",X"C6",
		X"6C",X"40",X"0C",X"60",X"00",X"00",X"00",X"94",X"46",X"0C",X"60",X"00",X"00",X"0C",X"0C",X"66",
		X"0C",X"70",X"00",X"00",X"70",X"00",X"68",X"57",X"70",X"00",X"00",X"00",X"00",X"68",X"59",X"50",
		X"00",X"00",X"00",X"00",X"68",X"45",X"40",X"00",X"00",X"00",X"06",X"68",X"44",X"40",X"00",X"00",
		X"00",X"0C",X"59",X"00",X"00",X"00",X"00",X"00",X"07",X"70",X"70",X"00",X"00",X"00",X"00",X"07",
		X"00",X"07",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"40",X"00",X"00",X"54",X"40",X"00",X"04",
		X"50",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"75",X"45",X"50",X"00",X"00",
		X"07",X"70",X"77",X"54",X"55",X"00",X"00",X"00",X"77",X"77",X"55",X"55",X"00",X"00",X"00",X"47",
		X"75",X"54",X"00",X"00",X"00",X"00",X"00",X"77",X"55",X"00",X"00",X"00",X"00",X"00",X"0D",X"DD",
		X"00",X"00",X"00",X"00",X"00",X"D6",X"66",X"C0",X"00",X"00",X"00",X"96",X"66",X"8C",X"6C",X"00",
		X"00",X"00",X"C6",X"6C",X"40",X"06",X"80",X"00",X"00",X"00",X"04",X"46",X"06",X"C0",X"00",X"00",
		X"00",X"06",X"67",X"6C",X"00",X"00",X"00",X"00",X"05",X"77",X"00",X"00",X"00",X"00",X"00",X"05",
		X"85",X"00",X"00",X"00",X"00",X"00",X"04",X"54",X"00",X"00",X"00",X"00",X"00",X"04",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",
		X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"07",X"40",X"00",X"00",X"00",X"00",X"00",
		X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"07",X"54",X"55",
		X"00",X"00",X"00",X"77",X"07",X"75",X"45",X"50",X"00",X"00",X"07",X"77",X"75",X"55",X"50",X"00",
		X"00",X"04",X"77",X"55",X"40",X"00",X"00",X"00",X"00",X"07",X"75",X"50",X"00",X"00",X"00",X"00",
		X"00",X"DD",X"D0",X"00",X"00",X"00",X"00",X"0D",X"66",X"00",X"00",X"00",X"00",X"09",X"66",X"C6",
		X"00",X"00",X"00",X"00",X"0C",X"6C",X"66",X"00",X"00",X"00",X"00",X"00",X"06",X"6C",X"00",X"00",
		X"00",X"00",X"00",X"66",X"CC",X"60",X"00",X"00",X"00",X"06",X"60",X"C6",X"60",X"00",X"00",X"00",
		X"77",X"00",X"66",X"60",X"00",X"00",X"00",X"49",X"40",X"66",X"66",X"00",X"00",X"00",X"45",X"40",
		X"70",X"06",X"00",X"00",X"00",X"44",X"49",X"00",X"07",X"70",X"00",X"00",X"00",X"07",X"00",X"00",
		X"70",X"00",X"00",X"00",X"75",X"00",X"00",X"07",X"40",X"00",X"07",X"05",X"00",X"00",X"00",X"40",
		X"00",X"45",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"44",X"00",X"00",X"00",X"00",
		X"05",X"77",X"77",X"75",X"00",X"00",X"00",X"57",X"AA",X"7A",X"A7",X"50",X"00",X"00",X"57",X"A7",
		X"77",X"A7",X"50",X"00",X"00",X"55",X"77",X"57",X"75",X"50",X"00",X"00",X"05",X"77",X"77",X"75",
		X"00",X"00",X"00",X"00",X"57",X"77",X"50",X"00",X"00",X"00",X"0D",X"DC",X"7C",X"DD",X"00",X"00",
		X"00",X"0C",X"CD",X"4D",X"CC",X"00",X"00",X"00",X"C6",X"6C",X"DC",X"66",X"C0",X"00",X"00",X"66",
		X"66",X"66",X"66",X"60",X"00",X"00",X"C6",X"C5",X"55",X"C6",X"C0",X"00",X"00",X"C9",X"75",X"85",
		X"79",X"C0",X"00",X"00",X"07",X"75",X"55",X"77",X"00",X"00",X"00",X"07",X"75",X"45",X"77",X"00",
		X"00",X"00",X"00",X"54",X"44",X"50",X"00",X"00",X"00",X"00",X"44",X"44",X"40",X"00",X"00",X"00",
		X"00",X"88",X"88",X"80",X"00",X"00",X"00",X"00",X"66",X"66",X"60",X"00",X"00",X"00",X"00",X"09",
		X"09",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"00",
		X"00",X"00",X"00",X"00",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"57",X"57",X"50",X"00",X"00",
		X"00",X"00",X"44",X"54",X"40",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"05",
		X"54",X"57",X"00",X"00",X"00",X"00",X"54",X"45",X"77",X"07",X"77",X"00",X"00",X"55",X"45",X"77",
		X"77",X"70",X"00",X"00",X"00",X"55",X"55",X"77",X"40",X"00",X"00",X"00",X"45",X"55",X"77",X"00",
		X"00",X"00",X"00",X"55",X"57",X"70",X"00",X"00",X"00",X"00",X"DD",X"DD",X"00",X"00",X"00",X"00",
		X"08",X"66",X"6D",X"D0",X"00",X"00",X"00",X"86",X"68",X"66",X"66",X"00",X"00",X"00",X"66",X"00",
		X"C6",X"66",X"60",X"00",X"06",X"60",X"00",X"4C",X"66",X"C0",X"00",X"06",X"60",X"C6",X"44",X"90",
		X"00",X"00",X"07",X"70",X"66",X"6C",X"0C",X"00",X"00",X"57",X"75",X"86",X"60",X"07",X"00",X"00",
		X"49",X"95",X"86",X"60",X"00",X"70",X"00",X"45",X"54",X"86",X"60",X"00",X"00",X"00",X"44",X"44",
		X"8C",X"60",X"00",X"00",X"00",X"44",X"44",X"8C",X"66",X"00",X"00",X"00",X"00",X"09",X"05",X"C0",
		X"00",X"00",X"00",X"00",X"07",X"07",X"70",X"00",X"00",X"00",X"00",X"70",X"00",X"70",X"00",X"00",
		X"00",X"54",X"00",X"00",X"07",X"00",X"00",X"00",X"05",X"00",X"00",X"04",X"70",X"00",X"00",X"05",
		X"50",X"00",X"04",X"04",X"40",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"05",X"54",
		X"57",X"00",X"00",X"00",X"00",X"54",X"45",X"77",X"07",X"77",X"00",X"00",X"55",X"45",X"77",X"77",
		X"70",X"00",X"00",X"00",X"55",X"55",X"77",X"40",X"00",X"00",X"00",X"45",X"55",X"77",X"00",X"00",
		X"00",X"00",X"55",X"57",X"70",X"00",X"00",X"00",X"00",X"DD",X"DD",X"00",X"00",X"00",X"00",X"00",
		X"C6",X"6D",X"D0",X"00",X"00",X"00",X"08",X"66",X"86",X"66",X"00",X"00",X"00",X"86",X"C0",X"C6",
		X"66",X"60",X"00",X"00",X"6C",X"00",X"4C",X"66",X"C0",X"00",X"00",X"C6",X"06",X"44",X"00",X"00",
		X"00",X"00",X"06",X"66",X"6C",X"00",X"00",X"00",X"00",X"00",X"77",X"60",X"00",X"00",X"00",X"00",
		X"00",X"77",X"50",X"00",X"00",X"00",X"00",X"05",X"88",X"50",X"00",X"00",X"00",X"00",X"04",X"55",
		X"40",X"00",X"00",X"00",X"00",X"04",X"44",X"40",X"00",X"00",X"00",X"00",X"04",X"44",X"40",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",
		X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"47",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"55",X"45",
		X"70",X"00",X"00",X"00",X"05",X"44",X"57",X"70",X"77",X"70",X"00",X"05",X"54",X"57",X"77",X"77",
		X"00",X"00",X"00",X"05",X"55",X"57",X"74",X"00",X"00",X"00",X"04",X"55",X"57",X"70",X"00",X"00",
		X"00",X"05",X"55",X"77",X"00",X"00",X"00",X"00",X"0D",X"DD",X"D0",X"00",X"00",X"00",X"00",X"00",
		X"66",X"DD",X"00",X"00",X"00",X"00",X"00",X"6C",X"66",X"60",X"00",X"00",X"00",X"00",X"6C",X"C6",
		X"66",X"00",X"00",X"00",X"00",X"66",X"C6",X"6C",X"00",X"00",X"00",X"00",X"C6",X"60",X"00",X"00",
		X"00",X"00",X"06",X"8C",X"66",X"00",X"00",X"00",X"00",X"06",X"C8",X"06",X"60",X"00",X"00",X"00",
		X"06",X"6C",X"00",X"77",X"00",X"00",X"00",X"06",X"66",X"00",X"77",X"50",X"00",X"00",X"66",X"6C",
		X"05",X"99",X"50",X"00",X"07",X"70",X"09",X"04",X"55",X"40",X"00",X"07",X"00",X"07",X"54",X"44",
		X"40",X"44",X"7E",X"00",X"00",X"04",X"44",X"40",X"04",X"70",X"00",X"00",X"50",X"00",X"00",X"54",
		X"00",X"00",X"00",X"04",X"70",X"00",X"40",X"00",X"00",X"00",X"04",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"05",X"50",X"00",X"00",X"05",X"50",X"00",X"00",X"00",X"00",X"05",X"55",X"55",X"50",
		X"00",X"00",X"00",X"45",X"55",X"4E",X"55",X"00",X"00",X"00",X"55",X"E5",X"4E",X"54",X"00",X"00",
		X"00",X"04",X"5E",X"E5",X"40",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"0D",
		X"DC",X"CD",X"D0",X"00",X"00",X"00",X"66",X"66",X"66",X"66",X"00",X"00",X"00",X"66",X"6C",X"C6",
		X"66",X"00",X"00",X"00",X"CC",X"94",X"49",X"CC",X"00",X"00",X"00",X"0E",X"9C",X"C9",X"E0",X"00",
		X"00",X"00",X"00",X"C6",X"6C",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"00",
		X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"70",X"00",X"00",X"00",X"00",X"00",X"07",X"70",X"00",
		X"00",X"00",X"00",X"00",X"07",X"70",X"00",X"00",X"00",X"00",X"00",X"E5",X"5E",X"00",X"00",X"00",
		X"00",X"00",X"5A",X"A5",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"05",
		X"54",X"57",X"00",X"00",X"00",X"00",X"55",X"45",X"77",X"07",X"70",X"00",X"00",X"55",X"55",X"77",
		X"77",X"00",X"00",X"00",X"00",X"45",X"57",X"74",X"00",X"00",X"00",X"00",X"55",X"77",X"00",X"00",
		X"00",X"00",X"00",X"DD",X"D0",X"00",X"00",X"00",X"00",X"06",X"66",X"6D",X"00",X"00",X"00",X"00",
		X"6C",X"08",X"66",X"69",X"00",X"00",X"06",X"C0",X"04",X"C6",X"6C",X"00",X"00",X"06",X"C0",X"64",
		X"49",X"00",X"00",X"00",X"07",X"C0",X"66",X"C0",X"C0",X"00",X"00",X"07",X"75",X"86",X"00",X"07",
		X"00",X"00",X"05",X"95",X"86",X"00",X"00",X"00",X"00",X"04",X"54",X"86",X"00",X"00",X"00",X"00",
		X"04",X"44",X"86",X"60",X"00",X"00",X"00",X"00",X"00",X"95",X"C0",X"00",X"00",X"00",X"00",X"07",
		X"07",X"70",X"00",X"00",X"00",X"00",X"70",X"00",X"70",X"00",X"00",X"00",X"04",X"00",X"00",X"07",
		X"00",X"00",X"00",X"05",X"40",X"00",X"04",X"45",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"00",X"05",X"54",X"57",X"00",X"00",X"00",X"00",X"55",X"45",X"77",X"07",X"70",X"00",X"00",
		X"55",X"55",X"77",X"77",X"00",X"00",X"00",X"00",X"45",X"57",X"74",X"00",X"00",X"00",X"00",X"55",
		X"77",X"00",X"00",X"00",X"00",X"00",X"DD",X"D0",X"00",X"00",X"00",X"00",X"0C",X"66",X"6D",X"00",
		X"00",X"00",X"00",X"C6",X"C8",X"66",X"69",X"00",X"00",X"08",X"60",X"04",X"C6",X"6C",X"00",X"00",
		X"0C",X"60",X"64",X"40",X"00",X"00",X"00",X"00",X"C6",X"76",X"60",X"00",X"00",X"00",X"00",X"00",
		X"77",X"50",X"00",X"00",X"00",X"00",X"00",X"58",X"50",X"00",X"00",X"00",X"00",X"00",X"45",X"40",
		X"00",X"00",X"00",X"00",X"00",X"44",X"40",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"70",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"00",X"00",X"55",X"45",X"70",X"00",X"00",X"00",X"05",X"54",X"57",X"70",
		X"77",X"00",X"00",X"05",X"55",X"57",X"77",X"70",X"00",X"00",X"00",X"04",X"55",X"77",X"40",X"00",
		X"00",X"00",X"05",X"57",X"70",X"00",X"00",X"00",X"00",X"0D",X"DD",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"D0",X"00",X"00",X"00",X"00",X"00",X"6C",X"66",X"90",X"00",X"00",X"00",X"00",X"66",
		X"C6",X"C0",X"00",X"00",X"00",X"00",X"C6",X"60",X"00",X"00",X"00",X"00",X"06",X"CC",X"66",X"00",
		X"00",X"00",X"00",X"06",X"6C",X"06",X"60",X"00",X"00",X"00",X"06",X"66",X"00",X"77",X"00",X"00",
		X"00",X"66",X"66",X"04",X"94",X"00",X"00",X"00",X"60",X"07",X"04",X"54",X"00",X"00",X"07",X"70",
		X"00",X"94",X"44",X"00",X"00",X"07",X"00",X"00",X"70",X"00",X"00",X"04",X"70",X"00",X"00",X"57",
		X"00",X"00",X"04",X"00",X"00",X"00",X"50",X"70",X"00",X"40",X"00",X"00",X"00",X"00",X"54",X"00",
		X"00",X"FE",X"4E",X"F0",X"00",X"00",X"0F",X"55",X"55",X"5F",X"00",X"00",X"F5",X"5E",X"4E",X"55",
		X"F0",X"00",X"0F",X"5E",X"EE",X"5F",X"00",X"00",X"00",X"FE",X"EE",X"F0",X"00",X"00",X"00",X"F6",
		X"66",X"F0",X"00",X"00",X"0F",X"66",X"66",X"6F",X"00",X"00",X"0F",X"C6",X"46",X"CF",X"00",X"00",
		X"0F",X"E5",X"45",X"EF",X"00",X"00",X"00",X"F6",X"66",X"F0",X"00",X"00",X"00",X"F6",X"66",X"F0",
		X"00",X"00",X"00",X"F6",X"66",X"F0",X"00",X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"00",X"0F",
		X"7F",X"00",X"00",X"00",X"00",X"0F",X"4F",X"00",X"00",X"00",X"00",X"F5",X"55",X"F0",X"00",X"00",
		X"00",X"0F",X"45",X"FF",X"00",X"00",X"0F",X"FF",X"74",X"55",X"F0",X"00",X"F7",X"7F",X"75",X"45",
		X"F0",X"00",X"0F",X"47",X"75",X"5F",X"00",X"00",X"00",X"FF",X"75",X"5F",X"00",X"00",X"00",X"0F",
		X"FD",X"D8",X"F0",X"00",X"00",X"FC",X"D6",X"66",X"6F",X"00",X"00",X"F6",X"64",X"00",X"C6",X"F0",
		X"00",X"0F",X"F4",X"6C",X"06",X"F0",X"00",X"00",X"FC",X"66",X"07",X"F0",X"00",X"07",X"FF",X"68",
		X"57",X"F0",X"00",X"00",X"F6",X"68",X"44",X"F0",X"00",X"00",X"0F",X"CF",X"44",X"F0",X"00",X"00",
		X"F7",X"F7",X"FF",X"00",X"00",X"FF",X"7F",X"0F",X"7F",X"00",X"0F",X"44",X"5F",X"0F",X"55",X"F0",
		X"00",X"0F",X"45",X"FF",X"00",X"00",X"0F",X"FF",X"74",X"55",X"F0",X"00",X"F7",X"7F",X"75",X"45",
		X"F0",X"00",X"0F",X"47",X"75",X"5F",X"00",X"00",X"00",X"FF",X"75",X"5F",X"00",X"00",X"00",X"0F",
		X"FD",X"D8",X"F0",X"00",X"00",X"FC",X"D6",X"66",X"8F",X"00",X"00",X"F6",X"64",X"FF",X"6F",X"00",
		X"00",X"0F",X"F4",X"68",X"6F",X"00",X"00",X"00",X"F6",X"67",X"F0",X"00",X"00",X"00",X"F5",X"77",
		X"F0",X"00",X"00",X"00",X"F5",X"5F",X"00",X"00",X"00",X"00",X"F4",X"4F",X"00",X"00",X"00",X"00",
		X"0F",X"7F",X"00",X"00",X"00",X"00",X"0F",X"7F",X"00",X"00",X"00",X"00",X"F4",X"4F",X"00",X"00",
		X"00",X"F4",X"5F",X"F0",X"00",X"00",X"FF",X"F7",X"45",X"5F",X"00",X"00",X"77",X"F7",X"54",X"5F",
		X"00",X"00",X"F4",X"77",X"55",X"F0",X"00",X"00",X"0F",X"F7",X"55",X"F0",X"00",X"00",X"00",X"FF",
		X"DD",X"F0",X"00",X"00",X"0F",X"CD",X"6F",X"00",X"00",X"00",X"0F",X"6C",X"6F",X"00",X"00",X"00",
		X"00",X"FF",X"66",X"F0",X"00",X"00",X"00",X"F6",X"C6",X"F0",X"00",X"00",X"0F",X"7F",X"66",X"F0",
		X"00",X"00",X"F4",X"4F",X"66",X"6F",X"00",X"00",X"F4",X"4F",X"FF",X"7F",X"00",X"00",X"0F",X"F7",
		X"F0",X"F7",X"F0",X"00",X"0F",X"7F",X"00",X"0F",X"4F",X"00",X"F5",X"5F",X"00",X"00",X"F4",X"00",
		X"00",X"FE",X"4E",X"F0",X"00",X"00",X"0F",X"57",X"77",X"5F",X"00",X"00",X"F5",X"50",X"70",X"55",
		X"F0",X"00",X"0F",X"57",X"77",X"5F",X"00",X"00",X"00",X"F5",X"75",X"F0",X"00",X"00",X"00",X"FD",
		X"4D",X"F0",X"00",X"00",X"0F",X"66",X"D6",X"6F",X"00",X"00",X"0F",X"C6",X"66",X"CF",X"00",X"00",
		X"0F",X"75",X"55",X"7F",X"00",X"00",X"00",X"F5",X"85",X"F0",X"00",X"00",X"00",X"F4",X"44",X"F0",
		X"00",X"00",X"00",X"F6",X"66",X"F0",X"00",X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"00",X"0F",
		X"7F",X"00",X"00",X"00",X"00",X"0F",X"7F",X"00",X"00",X"00",X"00",X"F4",X"54",X"F0",X"00",X"00",
		X"00",X"0F",X"F5",X"4F",X"00",X"00",X"00",X"F5",X"54",X"7F",X"FF",X"00",X"00",X"F5",X"45",X"7F",
		X"77",X"F0",X"00",X"0F",X"55",X"77",X"4F",X"00",X"00",X"0F",X"55",X"7F",X"F0",X"00",X"00",X"F8",
		X"DD",X"FF",X"00",X"00",X"0F",X"66",X"66",X"DC",X"F0",X"00",X"F6",X"C0",X"04",X"66",X"F0",X"00",
		X"F6",X"0C",X"64",X"FF",X"00",X"00",X"F7",X"06",X"6F",X"F0",X"00",X"00",X"F7",X"58",X"6F",X"F7",
		X"00",X"00",X"F4",X"48",X"66",X"F0",X"00",X"00",X"F4",X"4F",X"CF",X"00",X"00",X"00",X"0F",X"F7",
		X"F7",X"F0",X"00",X"00",X"0F",X"7F",X"0F",X"7F",X"F0",X"00",X"F5",X"5F",X"0F",X"54",X"4F",X"00",
		X"00",X"FF",X"54",X"F0",X"00",X"00",X"0F",X"55",X"47",X"FF",X"F0",X"00",X"0F",X"54",X"57",X"F7",
		X"7F",X"00",X"00",X"F5",X"57",X"74",X"F0",X"00",X"00",X"F5",X"57",X"FF",X"00",X"00",X"0F",X"8D",
		X"DF",X"F0",X"00",X"00",X"F8",X"66",X"6D",X"CF",X"00",X"00",X"F6",X"FF",X"46",X"6F",X"00",X"00",
		X"F6",X"86",X"4F",X"F0",X"F0",X"00",X"0F",X"76",X"6F",X"00",X"00",X"00",X"0F",X"77",X"5F",X"00",
		X"00",X"00",X"00",X"F5",X"5F",X"00",X"00",X"00",X"00",X"F4",X"4F",X"00",X"00",X"00",X"00",X"F7",
		X"F0",X"00",X"00",X"00",X"00",X"F7",X"F0",X"00",X"00",X"00",X"00",X"F4",X"4F",X"00",X"00",X"00",
		X"00",X"0F",X"F5",X"4F",X"00",X"00",X"00",X"F5",X"54",X"7F",X"FF",X"00",X"00",X"F5",X"45",X"7F",
		X"77",X"00",X"00",X"0F",X"55",X"77",X"4F",X"00",X"00",X"0F",X"55",X"7F",X"F0",X"00",X"00",X"0F",
		X"DD",X"FF",X"00",X"00",X"00",X"00",X"F6",X"DC",X"F0",X"00",X"00",X"00",X"F6",X"C6",X"F0",X"00",
		X"00",X"0F",X"66",X"FF",X"00",X"00",X"00",X"0F",X"6C",X"6F",X"00",X"00",X"00",X"0F",X"66",X"F7",
		X"F0",X"00",X"00",X"F6",X"66",X"F4",X"4F",X"00",X"00",X"F7",X"FF",X"F4",X"4F",X"00",X"0F",X"7F",
		X"0F",X"7F",X"F0",X"00",X"F4",X"F0",X"00",X"F7",X"F0",X"00",X"4F",X"00",X"00",X"F5",X"5F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"90",X"00",
		X"86",X"6C",X"CC",X"80",X"08",X"89",X"99",X"00",X"66",X"68",X"88",X"80",X"06",X"86",X"98",X"00",
		X"06",X"86",X"98",X"00",X"06",X"86",X"A8",X"00",X"06",X"86",X"A8",X"00",X"06",X"A6",X"A8",X"00",
		X"06",X"96",X"98",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"50",X"06",X"80",X"00",X"00",X"00",X"60",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"88",X"60",X"04",X"E0",X"06",X"00",X"B0",X"00",X"00",X"00",X"EB",
		X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"0B",X"B4",X"00",X"00",X"60",X"00",X"00",X"E4",X"2D",
		X"B0",X"00",X"06",X"00",X"86",X"00",X"00",X"42",X"00",X"06",X"68",X"00",X"08",X"60",X"00",X"52",
		X"00",X"00",X"80",X"00",X"00",X"80",X"05",X"0B",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"04",
		X"0B",X"50",X"00",X"00",X"00",X"06",X"00",X"40",X"00",X"00",X"60",X"00",X"00",X"86",X"00",X"50",
		X"00",X"00",X"60",X"00",X"00",X"00",X"05",X"00",X"06",X"00",X"00",X"00",X"00",X"40",X"00",X"00",
		X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"68",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"B0",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",
		X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"BF",X"B0",X"B0",X"00",X"00",X"00",X"0B",X"B4",
		X"44",X"4F",X"44",X"BB",X"00",X"00",X"00",X"0B",X"45",X"F4",X"4E",X"F4",X"44",X"00",X"00",X"00",
		X"B4",X"40",X"E0",X"FB",X"05",X"F4",X"B0",X"00",X"0B",X"44",X"40",X"BB",X"BE",X"5F",X"B0",X"5B",
		X"00",X"0B",X"45",X"5F",X"BE",X"4B",X"F0",X"4B",X"04",X"00",X"04",X"FF",X"0F",X"F0",X"5F",X"0B",
		X"44",X"BF",X"00",X"B4",X"E0",X"BA",X"5B",X"54",X"E4",X"F0",X"BB",X"00",X"44",X"FB",X"40",X"BF",
		X"44",X"EF",X"E4",X"44",X"00",X"4F",X"0B",X"04",X"05",X"EF",X"E0",X"0E",X"4F",X"00",X"00",X"00",
		X"0E",X"EF",X"EE",X"FE",X"00",X"00",X"00",X"00",X"00",X"4F",X"0F",X"5E",X"FF",X"BB",X"00",X"00",
		X"00",X"0B",X"40",X"0F",X"5F",X"00",X"FB",X"B0",X"00",X"00",X"04",X"F0",X"FE",X"EF",X"00",X"44",
		X"40",X"00",X"00",X"00",X"00",X"FE",X"EF",X"00",X"F4",X"F0",X"00",X"00",X"00",X"00",X"0A",X"E5",
		X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"0F",X"E5",X"00",X"00",X"00",X"00",X"00",X"00",X"07",
		X"07",X"57",X"07",X"00",X"00",X"00",X"00",X"00",X"07",X"77",X"77",X"77",X"00",X"00",X"00",X"00",
		X"00",X"07",X"F7",X"E7",X"F7",X"00",X"00",X"00",X"00",X"00",X"07",X"F7",X"E7",X"F7",X"00",X"00",
		X"00",X"00",X"00",X"07",X"F7",X"E7",X"A7",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"EF",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",
		X"0F",X"E0",X"00",X"00",X"00",X"00",X"0E",X"05",X"0F",X"5E",X"F0",X"50",X"00",X"00",X"00",X"50",
		X"50",X"E0",X"FE",X"0B",X"F0",X"00",X"00",X"00",X"0E",X"F0",X"40",X"BE",X"54",X"50",X"50",X"00",
		X"00",X"EB",X"54",X"4E",X"FB",X"F4",X"0E",X"00",X"00",X"0E",X"00",X"04",X"40",X"5F",X"00",X"EB",
		X"04",X"00",X"00",X"E4",X"E4",X"4F",X"54",X"EB",X"FB",X"0E",X"00",X"E0",X"44",X"40",X"BF",X"B4",
		X"EF",X"40",X"E0",X"00",X"0B",X"4B",X"40",X"05",X"EF",X"40",X"0E",X"00",X"00",X"40",X"40",X"4E",
		X"EB",X"EB",X"FE",X"0B",X"04",X"00",X"40",X"40",X"0B",X"4F",X"5E",X"F0",X"4B",X"04",X"00",X"40",
		X"00",X"B0",X"44",X"5F",X"00",X"44",X"00",X"00",X"04",X"04",X"00",X"FE",X"EF",X"40",X"B0",X"B0",
		X"00",X"04",X"04",X"00",X"F4",X"EF",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"0A",X"EB",X"F0",
		X"B0",X"40",X"00",X"04",X"00",X"00",X"0F",X"E5",X"F0",X"00",X"B0",X"00",X"00",X"00",X"07",X"07",
		X"57",X"F7",X"00",X"00",X"00",X"00",X"00",X"07",X"77",X"77",X"77",X"00",X"04",X"00",X"00",X"00",
		X"07",X"F7",X"E7",X"F7",X"00",X"00",X"00",X"00",X"00",X"07",X"F7",X"E7",X"F7",X"00",X"00",X"00",
		X"00",X"00",X"07",X"F7",X"E7",X"A7",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"50",X"EF",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"0F",
		X"E0",X"00",X"00",X"00",X"00",X"0E",X"05",X"0F",X"5E",X"F0",X"50",X"00",X"00",X"00",X"50",X"50",
		X"E0",X"FE",X"05",X"F0",X"00",X"00",X"00",X"0E",X"F0",X"E0",X"FE",X"5F",X"50",X"50",X"00",X"00",
		X"E5",X"5F",X"0E",X"F5",X"F0",X"0E",X"00",X"00",X"0E",X"00",X"0F",X"F0",X"5F",X"00",X"EF",X"00",
		X"00",X"00",X"E0",X"EA",X"5F",X"5F",X"EE",X"F0",X"0E",X"00",X"E0",X"00",X"00",X"EF",X"EE",X"EF",
		X"E0",X"E0",X"00",X"00",X"00",X"00",X"05",X"EF",X"E0",X"0E",X"00",X"00",X"00",X"00",X"0E",X"EF",
		X"EE",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"5E",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"5F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"EF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"E5",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"E5",X"F0",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"57",
		X"F7",X"00",X"00",X"00",X"00",X"00",X"07",X"77",X"77",X"77",X"00",X"00",X"00",X"00",X"0B",X"47",
		X"F7",X"E7",X"F7",X"4B",X"00",X"00",X"0B",X"44",X"B7",X"B7",X"B7",X"4B",X"4B",X"B0",X"00",X"44",
		X"B4",X"07",X"44",X"B7",X"4B",X"44",X"B4",X"00",X"00",X"04",X"40",X"44",X"47",X"00",X"44",X"00",
		X"00",X"00",X"00",X"B4",X"00",X"00",X"00",X"0B",X"4B",X"4E",X"B0",X"00",X"00",X"4E",X"FB",X"FE",
		X"4B",X"40",X"00",X"04",X"BF",X"0E",X"0E",X"40",X"00",X"4B",X"05",X"44",X"E0",X"F4",X"00",X"40",
		X"EE",X"BB",X"54",X"44",X"00",X"04",X"00",X"54",X"4E",X"40",X"00",X"BB",X"4B",X"E4",X"EF",X"FB",
		X"00",X"40",X"44",X"EE",X"FB",X"44",X"00",X"0E",X"40",X"FE",X"FB",X"40",X"00",X"0F",X"0F",X"EF",
		X"00",X"40",X"00",X"00",X"0F",X"5E",X"F0",X"00",X"00",X"00",X"00",X"F5",X"F0",X"00",X"00",X"00",
		X"00",X"FE",X"F0",X"00",X"00",X"00",X"0F",X"77",X"F0",X"00",X"00",X"00",X"0F",X"77",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"FE",X"00",X"00",X"00",X"0E",X"F0",X"FE",
		X"00",X"00",X"00",X"00",X"EF",X"0E",X"0E",X"00",X"00",X"00",X"45",X"0F",X"E0",X"FE",X"00",X"00",
		X"4E",X"44",X"54",X"E0",X"00",X"B0",X"00",X"5F",X"5E",X"00",X"00",X"4E",X"FE",X"B4",X"E4",X"BE",
		X"00",X"00",X"4F",X"EB",X"FE",X"44",X"00",X"0E",X"F0",X"4E",X"F4",X"04",X"00",X"0B",X"4F",X"B4",
		X"B0",X"40",X"00",X"4B",X"0F",X"5E",X"FB",X"0B",X"00",X"00",X"40",X"F5",X"F4",X"00",X"00",X"04",
		X"00",X"FE",X"F0",X"04",X"00",X"00",X"0F",X"77",X"F0",X"00",X"00",X"00",X"0F",X"77",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"FE",X"00",X"00",X"00",X"0E",X"F0",X"FE",
		X"00",X"00",X"00",X"00",X"EF",X"0E",X"0E",X"00",X"00",X"00",X"05",X"0F",X"E0",X"FE",X"00",X"00",
		X"EE",X"FF",X"5F",X"E0",X"00",X"00",X"00",X"5F",X"5E",X"00",X"00",X"EE",X"FE",X"5F",X"EF",X"FE",
		X"00",X"00",X"EF",X"EE",X"FE",X"EF",X"00",X"0E",X"F0",X"FE",X"F0",X"00",X"00",X"0F",X"0F",X"EF",
		X"00",X"00",X"00",X"00",X"0F",X"5E",X"F0",X"00",X"00",X"00",X"00",X"F5",X"F0",X"00",X"00",X"00",
		X"00",X"FE",X"F0",X"00",X"00",X"00",X"0F",X"77",X"F0",X"00",X"00",X"4B",X"0B",X"4E",X"B4",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"50",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E5",X"00",X"00",X"40",X"04",X"00",X"00",X"05",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"40",X"00",X"40",X"04",X"00",X"40",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"04",X"40",X"42",X"00",X"40",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"04",X"44",X"42",X"44",X"44",X"44",X"40",X"00",X"00",X"00",X"00",X"45",X"00",X"04",X"04",
		X"24",X"24",X"22",X"42",X"44",X"24",X"00",X"00",X"5E",X"00",X"00",X"04",X"44",X"04",X"42",X"44",
		X"24",X"42",X"22",X"42",X"44",X"40",X"44",X"00",X"00",X"00",X"00",X"04",X"44",X"24",X"D4",X"22",
		X"DD",X"24",X"22",X"44",X"44",X"40",X"00",X"00",X"00",X"00",X"04",X"24",X"44",X"2D",X"2D",X"D2",
		X"D2",X"D2",X"44",X"40",X"00",X"00",X"00",X"00",X"00",X"04",X"42",X"D2",X"42",X"D2",X"DD",X"DD",
		X"24",X"42",X"44",X"40",X"00",X"00",X"E5",X"40",X"44",X"44",X"4D",X"2D",X"DD",X"DD",X"DD",X"D2",
		X"D2",X"22",X"24",X"45",X"00",X"00",X"04",X"22",X"2D",X"22",X"DD",X"DD",X"DD",X"D2",X"22",X"44",
		X"40",X"00",X"00",X"00",X"00",X"00",X"44",X"44",X"42",X"2D",X"D2",X"22",X"D2",X"44",X"42",X"44",
		X"00",X"00",X"00",X"00",X"00",X"44",X"24",X"24",X"4D",X"22",X"42",X"2D",X"22",X"44",X"00",X"00",
		X"00",X"00",X"00",X"04",X"44",X"42",X"24",X"22",X"42",X"4D",X"44",X"44",X"20",X"00",X"00",X"00",
		X"00",X"00",X"45",X"00",X"04",X"44",X"44",X"24",X"42",X"42",X"40",X"44",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"00",X"40",X"00",X"02",X"40",X"44",X"00",X"40",X"00",X"00",X"00",X"00",
		X"00",X"04",X"44",X"00",X"40",X"00",X"04",X"40",X"04",X"00",X"54",X"E0",X"00",X"00",X"00",X"00",
		X"04",X"00",X"00",X"45",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",
		X"00",X"00",X"04",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0D",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"0D",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"BC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"5B",X"45",X"E0",X"0E",X"45",X"00",X"00",X"00",
		X"00",X"D0",X"00",X"00",X"E5",X"B4",X"B4",X"5E",X"5B",X"44",X"EE",X"00",X"00",X"00",X"06",X"00",
		X"00",X"0E",X"4B",X"45",X"5E",X"54",X"B4",X"45",X"E0",X"00",X"0D",X"60",X"00",X"00",X"55",X"55",
		X"4B",X"45",X"E5",X"4B",X"55",X"E5",X"E0",X"00",X"00",X"00",X"00",X"00",X"BB",X"44",X"55",X"5E",
		X"E4",X"45",X"5E",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",X"B5",X"5B",X"45",X"5E",X"54",X"B5",
		X"EE",X"EE",X"EE",X"00",X"D0",X"00",X"00",X"0E",X"44",X"E5",X"54",X"EE",X"E5",X"55",X"EE",X"EE",
		X"EE",X"00",X"60",X"00",X"D0",X"05",X"EB",X"4E",X"55",X"4E",X"5E",X"55",X"5E",X"EE",X"5E",X"00",
		X"00",X"00",X"D0",X"04",X"5E",X"45",X"EE",X"5E",X"55",X"EE",X"EE",X"E5",X"E0",X"00",X"00",X"00",
		X"00",X"0E",X"55",X"55",X"5E",X"E5",X"55",X"EE",X"55",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"55",X"EE",X"EE",X"EE",X"E5",X"EE",X"E0",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"0E",
		X"EE",X"EE",X"EE",X"EE",X"E0",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"D0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"00",X"00",X"D0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"0C",X"90",X"00",X"00",X"00",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EB",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E5",X"B4",X"5E",X"00",X"E4",X"50",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"5B",X"4B",X"45",X"E5",X"B4",X"4E",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E4",X"B4",X"55",X"E5",X"4B",X"44",
		X"5E",X"00",X"00",X"00",X"00",X"00",X"9C",X"00",X"00",X"00",X"05",X"55",X"54",X"B4",X"5E",X"54",
		X"B5",X"5E",X"5E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"0B",X"B4",X"45",X"55",
		X"EE",X"44",X"55",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"55",
		X"B4",X"55",X"E5",X"4B",X"5E",X"EE",X"EE",X"E0",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"E4",X"4E",X"55",X"4E",X"EE",X"55",X"5E",X"EE",X"EE",X"E0",X"00",X"00",X"09",X"00",X"00",X"00",
		X"00",X"00",X"5E",X"B4",X"E5",X"54",X"E5",X"E5",X"55",X"EE",X"E5",X"E0",X"00",X"00",X"00",X"00",
		X"0C",X"00",X"00",X"00",X"45",X"E4",X"5E",X"E5",X"E5",X"5E",X"EE",X"EE",X"5E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E5",X"55",X"55",X"EE",X"55",X"5E",X"E5",X"5E",X"E0",X"00",
		X"00",X"0C",X"C0",X"00",X"00",X"00",X"00",X"00",X"0E",X"E5",X"5E",X"EE",X"EE",X"EE",X"5E",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"C9",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E6",X"C0",X"00",X"00",X"00",X"00",
		X"E5",X"DD",X"5E",X"00",X"EC",X"60",X"00",X"00",X"00",X"0E",X"5B",X"CD",X"45",X"C5",X"B4",X"66",
		X"E0",X"00",X"00",X"00",X"E4",X"DD",X"55",X"65",X"4B",X"46",X"CE",X"00",X"00",X"05",X"55",X"56",
		X"B4",X"6E",X"5C",X"B5",X"DC",X"5E",X"00",X"00",X"06",X"D6",X"45",X"65",X"EC",X"44",X"56",X"CE",
		X"EE",X"00",X"00",X"06",X"C5",X"64",X"56",X"E5",X"4D",X"DC",X"EE",X"CE",X"E0",X"00",X"E4",X"CE",
		X"5D",X"4E",X"CE",X"56",X"CE",X"E6",X"6C",X"E0",X"00",X"5E",X"BD",X"E5",X"64",X"E5",X"E5",X"CC",
		X"DC",X"EC",X"E0",X"00",X"46",X"E4",X"DE",X"EC",X"E5",X"5E",X"CC",X"CC",X"CE",X"00",X"00",X"E5",
		X"DC",X"5C",X"EE",X"C5",X"5E",X"E5",X"CC",X"E0",X"00",X"00",X"0E",X"E5",X"CC",X"EE",X"EE",X"EC",
		X"CC",X"CE",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"6C",X"CC",X"EE",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"6C",X"00",X"00",X"00",X"00",X"00",X"0D",X"D0",X"00",X"00",X"C6",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"D0",X"0C",X"00",X"06",X"60",X"00",X"00",X"00",X"00",X"0D",X"D0",
		X"06",X"00",X"00",X"6C",X"00",X"00",X"00",X"00",X"00",X"60",X"06",X"00",X"C0",X"0D",X"C0",X"00",
		X"00",X"00",X"6D",X"60",X"06",X"00",X"C0",X"00",X"6C",X"00",X"00",X"00",X"00",X"6C",X"06",X"00",
		X"60",X"00",X"DD",X"C0",X"0C",X"00",X"00",X"00",X"0C",X"00",X"D0",X"0C",X"00",X"6C",X"00",X"66",
		X"C0",X"00",X"00",X"00",X"D0",X"06",X"00",X"00",X"0C",X"CD",X"C0",X"C0",X"00",X"00",X"60",X"0D",
		X"00",X"C0",X"00",X"0C",X"CC",X"C9",X"00",X"00",X"00",X"0D",X"C0",X"C0",X"0C",X"00",X"00",X"0C",
		X"C0",X"00",X"00",X"00",X"00",X"0C",X"CC",X"00",X"00",X"C9",X"C9",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C9",X"C9",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"04",X"00",
		X"50",X"00",X"00",X"00",X"00",X"00",X"50",X"04",X"05",X"00",X"00",X"00",X"00",X"04",X"00",X"04",
		X"22",X"4E",X"00",X"E5",X"00",X"05",X"00",X"24",X"42",X"2D",X"44",X"54",X"4E",X"00",X"00",X"54",
		X"22",X"42",X"D2",X"B2",X"24",X"50",X"00",X"05",X"B2",X"4D",X"2D",X"D2",X"D4",X"45",X"55",X"50",
		X"04",X"44",X"22",X"DD",X"DD",X"22",X"D2",X"44",X"00",X"04",X"22",X"2D",X"DD",X"DD",X"DD",X"24",
		X"25",X"00",X"44",X"4D",X"D2",X"2D",X"DD",X"D2",X"45",X"40",X"00",X"05",X"54",X"42",X"D2",X"D2",
		X"24",X"24",X"00",X"00",X"04",X"55",X"24",X"24",X"2D",X"44",X"50",X"40",X"00",X"00",X"00",X"45",
		X"45",X"24",X"20",X"05",X"00",X"00",X"00",X"05",X"00",X"05",X"55",X"04",X"00",X"00",X"00",X"00",
		X"00",X"05",X"05",X"05",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"0D",X"00",X"00",X"0D",X"00",X"00",
		X"E5",X"5E",X"E0",X"0E",X"CC",X"00",X"00",X"00",X"0E",X"5B",X"B4",X"45",X"E5",X"45",X"E0",X"00",
		X"00",X"0E",X"E4",X"B4",X"55",X"EB",X"B4",X"5E",X"00",X"00",X"D0",X"5B",X"55",X"E5",X"5E",X"B4",
		X"55",X"EE",X"E0",X"00",X"00",X"5B",X"4B",X"E5",X"E4",X"45",X"5E",X"EE",X"E0",X"D0",X"00",X"44",
		X"55",X"4E",X"E5",X"B5",X"EE",X"E5",X"E0",X"00",X"00",X"45",X"BE",X"55",X"E5",X"55",X"EE",X"5E",
		X"00",X"00",X"D0",X"E5",X"54",X"EE",X"EE",X"EE",X"55",X"50",X"0D",X"00",X"00",X"0E",X"E5",X"EE",
		X"55",X"E5",X"5E",X"00",X"00",X"00",X"00",X"00",X"0E",X"EE",X"EE",X"EE",X"00",X"D0",X"00",X"00",
		X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",
		X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E5",X"5E",X"E0",X"0E",X"CC",X"00",X"00",
		X"C0",X"00",X"00",X"0E",X"5B",X"B4",X"45",X"E5",X"45",X"E0",X"00",X"00",X"00",X"00",X"0E",X"E4",
		X"B4",X"55",X"EB",X"B4",X"5E",X"00",X"00",X"00",X"00",X"00",X"5B",X"55",X"E5",X"5E",X"B4",X"55",
		X"EE",X"E0",X"00",X"C0",X"00",X"00",X"5B",X"4B",X"E5",X"E4",X"45",X"5E",X"EE",X"E0",X"00",X"00",
		X"00",X"00",X"44",X"55",X"4E",X"E5",X"B5",X"EE",X"E5",X"E0",X"00",X"00",X"00",X"00",X"45",X"BE",
		X"55",X"E5",X"55",X"EE",X"5E",X"00",X"00",X"00",X"00",X"00",X"E5",X"54",X"EE",X"EE",X"EE",X"55",
		X"50",X"00",X"00",X"00",X"A0",X"00",X"0E",X"E5",X"EE",X"55",X"E5",X"5E",X"00",X"00",X"0C",X"00",
		X"00",X"00",X"00",X"0E",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",
		X"00",X"00",X"00",X"00",X"E5",X"5E",X"E0",X"0E",X"6C",X"00",X"00",X"0E",X"5B",X"B4",X"45",X"E5",
		X"46",X"E0",X"00",X"0E",X"E4",X"B6",X"55",X"EB",X"B4",X"CE",X"00",X"00",X"5B",X"56",X"E5",X"6E",
		X"B4",X"56",X"EE",X"E0",X"00",X"5B",X"4B",X"65",X"C6",X"46",X"DE",X"EE",X"E0",X"00",X"D4",X"65",
		X"46",X"E6",X"CD",X"EE",X"EC",X"E0",X"00",X"C5",X"B6",X"56",X"E6",X"5C",X"EE",X"56",X"00",X"00",
		X"E6",X"56",X"E6",X"E6",X"EC",X"CD",X"C0",X"00",X"00",X"0E",X"D6",X"E6",X"5C",X"EC",X"6E",X"00",
		X"00",X"00",X"00",X"0E",X"DC",X"DC",X"DE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",
		X"0C",X"00",X"60",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"60",X"CD",X"06",X"D0",X"00",X"00",
		X"00",X"D0",X"C0",X"0D",X"06",X"CD",X"00",X"0C",X"00",X"00",X"C0",X"0D",X"06",X"06",X"0C",X"00",
		X"06",X"00",X"00",X"06",X"06",X"06",X"06",X"0C",X"CD",X"C0",X"00",X"00",X"00",X"D6",X"06",X"0C",
		X"0C",X"60",X"00",X"00",X"00",X"00",X"00",X"6C",X"6C",X"60",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"28",X"43",X"29",X"20",X"31",X"39",
		X"38",X"34",X"2C",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",
		X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"D0",X"00",X"50",
		X"40",X"50",X"0D",X"00",X"00",X"50",X"54",X"24",X"E5",X"40",X"00",X"00",X"04",X"D2",X"D2",X"2D",
		X"50",X"00",X"00",X"E4",X"2D",X"DD",X"D2",X"45",X"00",X"50",X"42",X"DD",X"DD",X"DD",X"24",X"00",
		X"04",X"DD",X"2D",X"DD",X"24",X"5E",X"00",X"0E",X"E4",X"D2",X"D2",X"D5",X"E0",X"00",X"00",X"4E",
		X"54",X"24",X"54",X"05",X"00",X"00",X"00",X"50",X"40",X"50",X"00",X"00",X"D0",X"00",X"00",X"50",
		X"00",X"0D",X"00",X"00",X"00",X"00",X"0D",X"00",X"0D",X"00",X"00",X"D0",X"C0",X"0E",X"EE",X"40",
		X"00",X"0C",X"0E",X"44",X"54",X"B4",X"E0",X"00",X"00",X"EB",X"45",X"B4",X"5E",X"E0",X"C0",X"C0",
		X"B5",X"EE",X"45",X"EE",X"5E",X"00",X"0E",X"45",X"4E",X"55",X"EE",X"5E",X"00",X"DE",X"E5",X"E4",
		X"EE",X"55",X"E0",X"00",X"00",X"EE",X"EE",X"EE",X"E0",X"0D",X"00",X"00",X"0C",X"00",X"D0",X"C0",
		X"00",X"00",X"00",X"00",X"0A",X"00",X"09",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",
		X"D0",X"00",X"A0",X"00",X"00",X"00",X"EE",X"E4",X"00",X"00",X"00",X"00",X"E4",X"45",X"4B",X"4E",
		X"00",X"00",X"00",X"0E",X"B4",X"5B",X"45",X"EE",X"00",X"90",X"A0",X"0B",X"5E",X"E4",X"5E",X"E5",
		X"E0",X"00",X"00",X"E4",X"54",X"E5",X"5E",X"E5",X"E0",X"00",X"00",X"EE",X"5E",X"4E",X"E5",X"5E",
		X"00",X"00",X"90",X"0E",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"EE",X"E6",X"00",X"00",X"E4",
		X"4C",X"4B",X"CE",X"00",X"0E",X"B6",X"5B",X"C6",X"EE",X"00",X"06",X"5E",X"C4",X"DE",X"E5",X"E0",
		X"D4",X"64",X"65",X"CC",X"E6",X"E0",X"E6",X"CE",X"CE",X"E6",X"CE",X"00",X"0E",X"C6",X"D6",X"DE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",
		X"0C",X"00",X"C0",X"00",X"00",X"06",X"00",X"06",X"00",X"00",X"06",X"00",X"C0",X"D0",X"00",X"00",
		X"D0",X"60",X"60",X"CC",X"06",X"00",X"06",X"C0",X"C0",X"06",X"C0",X"00",X"00",X"C6",X"D6",X"D0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"EE",X"00",X"E4",X"E0",X"0E",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"45",X"EE",X"54",X"5E",
		X"E5",X"4E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"54",
		X"5E",X"52",X"5E",X"54",X"5E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E5",X"24",X"52",X"54",X"25",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"42",X"42",X"42",X"4E",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"55",X"54",X"23",X"24",X"55",X"5E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E4",X"42",X"22",X"33",X"32",X"22",
		X"44",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"55",X"54",
		X"23",X"24",X"55",X"5E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"42",X"42",X"42",X"4E",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E5",X"24",X"52",X"54",X"25",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"54",X"5E",X"52",X"5E",X"54",X"5E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"45",X"EE",X"54",X"5E",X"E5",X"4E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"EE",X"0E",X"54",
		X"5E",X"0E",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E4",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"40",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"04",X"20",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"04",
		X"00",X"02",X"00",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"02",X"40",X"00",X"20",X"02",X"40",X"02",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"44",X"40",X"44",X"00",X"44",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"44",X"02",X"42",X"40",X"40",X"42",X"00",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"00",X"42",X"24",X"44",X"42",X"44",X"42",
		X"24",X"44",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"42",X"24",
		X"42",X"24",X"22",X"42",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"00",X"42",X"22",X"42",X"22",X"22",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"04",X"02",X"44",X"42",X"22",X"22",X"22",X"44",X"40",X"40",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"42",X"22",X"23",X"22",X"22",X"44",X"24",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"42",X"22",X"22",X"22",X"33",X"32",X"22",X"22",
		X"20",X"22",X"42",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"22",X"22",X"22",X"23",
		X"22",X"22",X"42",X"40",X"04",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",
		X"42",X"22",X"22",X"22",X"22",X"44",X"42",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",
		X"00",X"00",X"42",X"42",X"22",X"22",X"22",X"24",X"42",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"44",X"22",X"24",X"22",X"24",X"22",X"24",X"40",X"00",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"04",X"24",X"24",X"42",X"44",X"44",X"22",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"44",X"04",X"22",X"44",
		X"04",X"42",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",
		X"40",X"22",X"44",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"04",X"00",X"00",X"42",X"40",X"00",X"00",X"02",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"24",X"00",X"04",X"00",X"40",X"00",X"00",X"00",X"44",X"20",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"20",X"20",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"40",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",
		X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"00",X"40",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"04",X"20",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"04",X"00",
		X"02",X"00",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"02",
		X"40",X"00",X"20",X"02",X"40",X"02",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"00",X"00",X"44",X"40",X"44",X"00",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"44",X"02",X"4F",X"40",X"40",X"42",X"00",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"00",X"42",X"24",X"44",X"4F",X"44",X"4F",X"F4",
		X"44",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"4F",X"F4",X"4F",
		X"F4",X"FF",X"42",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",
		X"4F",X"FF",X"4F",X"FF",X"FF",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",
		X"00",X"04",X"02",X"F4",X"4F",X"FF",X"FF",X"FF",X"44",X"40",X"40",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"24",X"4F",X"FF",X"FF",X"FF",X"FF",X"44",X"F4",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"4F",X"FF",X"FF",X"FF",X"F3",X"FF",X"FF",X"FF",X"F0",
		X"22",X"42",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"4F",X"40",X"04",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"4F",
		X"FF",X"FF",X"FF",X"FF",X"44",X"42",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",
		X"00",X"4F",X"4F",X"FF",X"FF",X"FF",X"F4",X"4F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"44",X"FF",X"FF",X"FF",X"F4",X"FF",X"F4",X"40",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"04",X"F4",X"F4",X"4F",X"4F",X"44",X"FF",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"44",X"04",X"FF",X"44",X"04",
		X"4F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"40",
		X"FF",X"44",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"04",X"00",X"00",X"4F",X"40",X"00",X"00",X"02",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"24",X"00",X"04",X"00",X"40",X"00",X"00",X"00",X"44",X"20",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"20",X"20",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"40",X"00",X"00",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"20",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"02",X"00",
		X"22",X"00",X"02",X"02",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"02",X"20",X"02",X"00",X"02",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"02",X"20",X"00",X"02",X"20",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"22",X"00",X"22",X"20",X"02",X"22",X"00",X"00",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"20",X"00",X"22",X"20",X"02",X"20",X"22",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"20",X"02",X"20",X"00",X"02",X"22",X"02",
		X"22",X"22",X"20",X"20",X"20",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"22",X"20",X"22",X"20",
		X"02",X"22",X"22",X"22",X"22",X"22",X"02",X"20",X"02",X"20",X"00",X"00",X"00",X"00",X"00",X"02",
		X"02",X"22",X"22",X"02",X"22",X"22",X"22",X"22",X"20",X"22",X"00",X"22",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"22",X"22",X"22",X"2F",X"22",X"20",X"22",X"22",X"22",X"20",X"00",
		X"00",X"00",X"00",X"00",X"22",X"20",X"22",X"02",X"22",X"22",X"22",X"2F",X"22",X"2F",X"F2",X"22",
		X"22",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"22",X"22",X"2F",X"F2",X"2F",X"F2",
		X"FF",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"22",X"2F",
		X"FF",X"2F",X"FF",X"FF",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"22",X"02",
		X"02",X"22",X"22",X"2F",X"FF",X"FF",X"FF",X"22",X"22",X"22",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"22",X"22",X"22",X"22",X"2F",X"FF",X"FF",X"FF",X"FF",X"22",X"F2",X"22",X"22",X"22",X"20",
		X"00",X"00",X"20",X"22",X"22",X"22",X"2F",X"FF",X"FF",X"FF",X"F3",X"FF",X"FF",X"FF",X"F0",X"22",
		X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"22",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"22",X"22",X"02",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"22",X"22",X"2F",X"FF",
		X"FF",X"FF",X"FF",X"22",X"22",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"22",
		X"2F",X"2F",X"FF",X"FF",X"FF",X"F2",X"2F",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"02",
		X"00",X"22",X"22",X"22",X"FF",X"FF",X"FF",X"F2",X"FF",X"F2",X"20",X"20",X"02",X"22",X"00",X"00",
		X"00",X"00",X"00",X"02",X"22",X"22",X"22",X"F2",X"F2",X"2F",X"2F",X"22",X"F2",X"22",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"22",X"20",X"00",X"22",X"22",X"02",X"FF",X"22",X"22",X"2F",
		X"22",X"22",X"20",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"22",X"22",X"22",X"FF",
		X"22",X"22",X"22",X"20",X"00",X"02",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"22",
		X"22",X"22",X"2F",X"22",X"22",X"22",X"22",X"20",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"22",X"00",X"22",X"22",X"22",X"20",X"22",X"20",X"22",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"20",X"02",X"22",X"22",X"22",X"20",X"22",X"00",X"22",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"22",X"02",X"22",X"22",X"20",X"02",X"20",X"00",
		X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"20",X"22",X"20",X"22",X"22",
		X"02",X"20",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"22",
		X"00",X"22",X"20",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"20",X"00",X"02",X"20",X"00",X"02",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"04",X"00",X"00",X"00",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"04",X"00",X"00",X"02",X"00",X"00",X"00",X"00",
		X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"04",X"40",X"04",
		X"20",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"02",X"00",X"02",
		X"00",X"40",X"00",X"20",X"40",X"04",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"04",X"02",X"40",X"00",X"04",X"00",X"04",X"00",X"00",X"00",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"40",X"00",X"24",X"04",X"04",X"20",X"44",X"00",X"00",
		X"24",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"04",X"42",X"00",X"20",
		X"40",X"04",X"02",X"44",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"20",X"04",X"00",X"00",
		X"02",X"00",X"04",X"00",X"40",X"20",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"04",X"02",X"00",
		X"04",X"40",X"00",X"40",X"00",X"00",X"00",X"02",X"04",X"00",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"00",X"04",X"40",X"00",X"44",X"44",X"00",X"00",X"DD",X"0F",X"DD",X"00",X"00",X"04",X"04",
		X"40",X"40",X"00",X"00",X"00",X"00",X"02",X"20",X"00",X"44",X"0C",X"DD",X"DC",X"CD",X"CC",X"DF",
		X"00",X"40",X"42",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"CC",X"D6",
		X"6D",X"CC",X"DD",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"20",X"02",X"00",X"00",X"40",
		X"0D",X"CC",X"CD",X"DC",X"CD",X"CC",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"00",X"40",X"00",X"00",X"DC",X"CC",X"CC",X"CC",X"66",X"6D",X"00",X"44",X"44",X"04",X"40",X"20",
		X"00",X"00",X"04",X"04",X"40",X"00",X"07",X"6C",X"76",X"CC",X"DD",X"6D",X"D0",X"00",X"22",X"00",
		X"00",X"00",X"00",X"00",X"04",X"40",X"00",X"00",X"00",X"07",X"6C",X"76",X"67",X"CC",X"DF",X"00",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"20",X"00",X"D6",X"67",X"7C",
		X"CC",X"DF",X"00",X"04",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"0D",X"DC",X"CD",X"CC",X"D0",X"0F",X"00",X"20",X"04",X"40",X"00",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"00",X"00",X"07",X"6C",X"6D",X"0F",X"40",X"04",X"02",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"20",X"00",X"40",X"07",X"66",X"D0",X"00",X"44",X"04",X"40",X"20",X"00",
		X"00",X"00",X"00",X"00",X"20",X"44",X"02",X"04",X"04",X"00",X"00",X"77",X"00",X"02",X"00",X"00",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"40",X"00",X"00",X"04",X"00",X"00",
		X"00",X"20",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"04",X"00",X"00",X"20",
		X"04",X"00",X"40",X"40",X"02",X"04",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",
		X"02",X"04",X"00",X"00",X"00",X"40",X"44",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"00",X"00",X"42",X"00",X"40",X"00",X"42",X"04",X"00",X"00",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"00",X"24",X"02",X"00",X"40",X"00",X"40",X"20",X"00",X"00",X"00",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"20",
		X"00",X"02",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"20",X"00",
		X"20",X"00",X"02",X"04",X"00",X"20",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"00",X"40",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DC",X"D0",X"00",X"00",X"0D",X"CC",
		X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"CC",X"CD",X"00",
		X"00",X"0C",X"CC",X"CD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DC",
		X"CC",X"CD",X"00",X"00",X"DC",X"CC",X"CD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0D",X"CC",X"CC",X"00",X"00",X"DC",X"CC",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"CC",X"00",X"00",X"CD",X"C0",X"00",X"0D",X"D0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",
		X"DC",X"CD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0D",X"CC",X"CD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"DC",X"DC",X"CC",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"DD",X"C0",X"00",X"00",X"00",X"00",X"00",X"DC",X"CD",X"CD",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0D",X"CC",X"CD",X"00",X"00",X"00",X"00",X"00",X"0D",X"D0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"CC",X"CD",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DC",X"D0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"CD",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"CD",X"CD",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DC",X"C0",X"00",X"00",X"00",X"0D",X"DC",X"CC",X"D0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"CC",X"C0",X"00",X"CC",X"00",X"00",
		X"DC",X"CC",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"CD",X"00",X"0D",
		X"CC",X"D0",X"00",X"DC",X"CD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"CC",
		X"CD",X"00",X"DC",X"CC",X"CD",X"00",X"0D",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0D",X"CC",X"D0",X"00",X"DC",X"DC",X"CD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"DD",X"00",X"00",X"DC",X"DC",X"CD",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"CD",X"D0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0D",X"CC",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"CC",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DC",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"D0",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"CD",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"CC",X"CD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"CC",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"0C",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"CC",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"D0",X"00",X"00",X"0C",X"CC",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"CC",X"D0",X"00",X"00",
		X"0D",X"CC",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"CC",
		X"D0",X"00",X"00",X"0D",X"CC",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"B0",X"BB",X"B0",X"BB",
		X"B0",X"BB",X"B0",X"00",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",X"BB",X"B0",X"B0",X"B0",X"B0",
		X"B0",X"B0",X"B0",X"B0",X"00",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",X"BB",X"B0",X"BB",X"B0",X"BB",
		X"B0",X"BB",X"B0",X"00",X"B0",X"BB",X"B0",X"BB",X"B0",X"BB",X"B0",X"00",X"B0",X"B0",X"B0",X"B0",
		X"B0",X"B0",X"B0",X"00",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",X"00",X"B0",X"B0",X"B0",X"B0",
		X"B0",X"B0",X"B0",X"00",X"B0",X"BB",X"B0",X"BB",X"B0",X"BB",X"B0",X"00",X"BB",X"B0",X"BB",X"B0",
		X"BB",X"B0",X"00",X"00",X"00",X"B0",X"B0",X"00",X"B0",X"B0",X"00",X"00",X"00",X"B0",X"BB",X"B0",
		X"B0",X"B0",X"00",X"00",X"00",X"B0",X"00",X"B0",X"B0",X"B0",X"00",X"00",X"00",X"B0",X"BB",X"B0",
		X"BB",X"B0",X"00",X"00",X"BB",X"B0",X"BB",X"B0",X"BB",X"B0",X"00",X"00",X"B0",X"00",X"B0",X"B0",
		X"B0",X"B0",X"00",X"00",X"BB",X"B0",X"B0",X"B0",X"B0",X"B0",X"00",X"00",X"00",X"B0",X"B0",X"B0",
		X"B0",X"B0",X"00",X"00",X"BB",X"B0",X"BB",X"B0",X"BB",X"B0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"11",X"11",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"11",X"11",X"00",X"11",X"00",X"11",X"00",
		X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",
		X"11",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"10",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"10",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",
		X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",
		X"11",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"28",X"43",X"29",X"20",X"31",X"39",
		X"38",X"34",X"2C",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",
		X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"60",X"33",X"00",
		X"67",X"6C",X"44",X"5C",X"45",X"72",X"72",X"6F",X"72",X"FF",X"60",X"40",X"00",X"5B",X"6C",X"66",
		X"5C",X"42",X"6F",X"78",X"20",X"6F",X"66",X"66",X"69",X"63",X"65",X"20",X"72",X"6F",X"62",X"62",
		X"65",X"72",X"79",X"21",X"5C",X"53",X"74",X"6F",X"70",X"20",X"74",X"68",X"65",X"20",X"68",X"65",
		X"69",X"73",X"74",X"21",X"FF",X"60",X"6B",X"00",X"64",X"6C",X"66",X"5C",X"47",X"75",X"61",X"72",
		X"64",X"20",X"61",X"67",X"61",X"69",X"6E",X"73",X"74",X"5C",X"6D",X"75",X"6C",X"74",X"69",X"70",
		X"6C",X"65",X"20",X"74",X"68",X"65",X"66",X"74",X"73",X"2E",X"FF",X"60",X"91",X"00",X"64",X"6C",
		X"66",X"5C",X"54",X"75",X"72",X"6B",X"65",X"79",X"20",X"61",X"69",X"72",X"20",X"72",X"61",X"69",
		X"64",X"21",X"5C",X"50",X"72",X"6F",X"74",X"65",X"63",X"74",X"20",X"74",X"68",X"65",X"5C",X"68",
		X"65",X"6C",X"69",X"63",X"6F",X"70",X"74",X"65",X"72",X"21",X"FF",X"60",X"C1",X"00",X"5E",X"6C",
		X"66",X"5C",X"41",X"6E",X"6F",X"6E",X"79",X"6D",X"6F",X"75",X"73",X"20",X"74",X"69",X"70",X"20",
		X"74",X"68",X"61",X"74",X"5C",X"48",X"69",X"2D",X"46",X"69",X"20",X"4E",X"6F",X"6F",X"6B",X"20",
		X"6D",X"61",X"79",X"20",X"62",X"65",X"5C",X"72",X"6F",X"62",X"62",X"65",X"64",X"2E",X"21",X"FF",
		X"60",X"F6",X"00",X"55",X"6C",X"66",X"5C",X"43",X"6C",X"6F",X"74",X"68",X"69",X"6E",X"67",X"20",
		X"73",X"74",X"6F",X"72",X"65",X"20",X"61",X"6C",X"61",X"72",X"6D",X"21",X"5C",X"44",X"65",X"73",
		X"69",X"67",X"6E",X"65",X"72",X"20",X"6A",X"65",X"61",X"6E",X"73",X"20",X"69",X"6E",X"5C",X"6A",
		X"65",X"6F",X"70",X"61",X"72",X"64",X"79",X"21",X"FF",X"61",X"2F",X"00",X"58",X"6C",X"66",X"5C",
		X"52",X"6F",X"62",X"62",X"65",X"72",X"79",X"20",X"69",X"6E",X"20",X"70",X"72",X"6F",X"67",X"72",
		X"65",X"73",X"73",X"21",X"5C",X"43",X"61",X"72",X"65",X"66",X"75",X"6C",X"21",X"5C",X"54",X"75",
		X"72",X"6B",X"65",X"79",X"73",X"20",X"64",X"69",X"73",X"67",X"75",X"69",X"73",X"65",X"64",X"20",
		X"61",X"73",X"5C",X"62",X"75",X"73",X"69",X"6E",X"65",X"73",X"73",X"6D",X"65",X"6E",X"21",X"FF",
		X"61",X"76",X"00",X"5E",X"6C",X"66",X"5C",X"4D",X"61",X"6A",X"6F",X"72",X"20",X"61",X"74",X"74",
		X"61",X"63",X"6B",X"20",X"69",X"73",X"5C",X"62",X"72",X"65",X"77",X"69",X"6E",X"67",X"21",X"20",
		X"20",X"50",X"72",X"6F",X"74",X"65",X"63",X"74",X"5C",X"74",X"68",X"65",X"20",X"68",X"65",X"6C",
		X"69",X"63",X"6F",X"70",X"74",X"65",X"72",X"20",X"61",X"6E",X"64",X"5C",X"61",X"6C",X"6C",X"20",
		X"73",X"74",X"6F",X"72",X"65",X"73",X"2E",X"FF",X"61",X"BE",X"00",X"55",X"6C",X"66",X"5C",X"54",
		X"75",X"72",X"6B",X"65",X"79",X"20",X"62",X"6F",X"6E",X"75",X"73",X"20",X"72",X"6F",X"75",X"6E",
		X"64",X"21",X"5C",X"54",X"65",X"72",X"6D",X"69",X"6E",X"61",X"74",X"65",X"20",X"61",X"73",X"20",
		X"6D",X"61",X"6E",X"79",X"5C",X"63",X"72",X"69",X"6D",X"69",X"6E",X"61",X"6C",X"73",X"20",X"61",
		X"73",X"20",X"70",X"6F",X"73",X"73",X"69",X"62",X"6C",X"65",X"5C",X"69",X"6E",X"20",X"31",X"35",
		X"20",X"73",X"65",X"63",X"6F",X"6E",X"64",X"73",X"2E",X"FF",X"62",X"16",X"00",X"73",X"9C",X"22",
		X"62",X"16",X"00",X"73",X"84",X"22",X"5C",X"52",X"61",X"70",X"69",X"64",X"20",X"46",X"69",X"72",
		X"65",X"21",X"FF",X"62",X"2F",X"00",X"5B",X"B4",X"22",X"62",X"2F",X"00",X"5B",X"9C",X"22",X"55",
		X"6E",X"6C",X"69",X"6D",X"69",X"74",X"65",X"64",X"20",X"47",X"72",X"65",X"6E",X"61",X"64",X"65",
		X"73",X"21",X"FF",X"62",X"49",X"00",X"5B",X"6C",X"66",X"5C",X"54",X"75",X"72",X"6B",X"65",X"79",
		X"20",X"62",X"6F",X"6E",X"75",X"73",X"20",X"72",X"6F",X"75",X"6E",X"64",X"21",X"FF",X"62",X"64",
		X"00",X"5B",X"6C",X"66",X"5C",X"54",X"75",X"72",X"6B",X"65",X"79",X"20",X"62",X"6C",X"69",X"74",
		X"7A",X"21",X"20",X"20",X"41",X"72",X"65",X"61",X"5C",X"75",X"6E",X"64",X"65",X"72",X"20",X"68",
		X"65",X"61",X"76",X"79",X"20",X"67",X"75",X"61",X"72",X"64",X"2E",X"FF",X"62",X"92",X"00",X"61",
		X"6C",X"66",X"5C",X"54",X"75",X"72",X"6B",X"65",X"79",X"20",X"61",X"69",X"72",X"20",X"72",X"61",
		X"69",X"64",X"21",X"5C",X"42",X"6C",X"61",X"73",X"74",X"20",X"74",X"68",X"65",X"6D",X"20",X"69",
		X"6E",X"20",X"74",X"68",X"65",X"5C",X"61",X"69",X"72",X"2E",X"FF",X"62",X"C1",X"00",X"58",X"6C",
		X"66",X"5C",X"43",X"79",X"62",X"6F",X"72",X"67",X"20",X"74",X"68",X"72",X"65",X"61",X"74",X"21",
		X"5C",X"54",X"75",X"72",X"6B",X"65",X"79",X"20",X"74",X"65",X"63",X"68",X"6E",X"6F",X"6C",X"6F",
		X"67",X"79",X"5C",X"77",X"69",X"6C",X"6C",X"20",X"61",X"74",X"74",X"65",X"6D",X"70",X"74",X"20",
		X"74",X"6F",X"5C",X"74",X"68",X"77",X"61",X"72",X"74",X"20",X"79",X"6F",X"75",X"72",X"20",X"65",
		X"66",X"66",X"6F",X"72",X"74",X"73",X"2E",X"FF",X"63",X"0E",X"00",X"67",X"6C",X"66",X"5C",X"53",
		X"68",X"6F",X"70",X"70",X"69",X"6E",X"67",X"20",X"73",X"70",X"72",X"65",X"65",X"21",X"5C",X"50",
		X"72",X"6F",X"74",X"65",X"63",X"74",X"20",X"74",X"68",X"65",X"5C",X"62",X"79",X"73",X"74",X"61",
		X"6E",X"64",X"65",X"72",X"73",X"2E",X"FF",X"63",X"3D",X"00",X"5E",X"6C",X"66",X"5C",X"4D",X"61",
		X"6A",X"6F",X"72",X"20",X"61",X"74",X"74",X"61",X"63",X"6B",X"20",X"69",X"73",X"5C",X"62",X"72",
		X"65",X"77",X"69",X"6E",X"67",X"21",X"20",X"20",X"50",X"72",X"6F",X"74",X"65",X"63",X"74",X"5C",
		X"61",X"6C",X"6C",X"20",X"6C",X"6F",X"63",X"61",X"74",X"69",X"6F",X"6E",X"73",X"20",X"66",X"72",
		X"6F",X"6D",X"5C",X"67",X"72",X"6F",X"75",X"6E",X"64",X"20",X"61",X"6E",X"64",X"20",X"61",X"69",
		X"72",X"5C",X"61",X"74",X"74",X"61",X"63",X"6B",X"21",X"FF",X"63",X"90",X"00",X"61",X"6C",X"66",
		X"5C",X"4C",X"61",X"73",X"74",X"20",X"73",X"74",X"61",X"6E",X"64",X"20",X"6F",X"66",X"20",X"74",
		X"68",X"65",X"5C",X"74",X"75",X"72",X"6B",X"65",X"79",X"73",X"2E",X"FF",X"63",X"B2",X"00",X"55",
		X"6C",X"66",X"5C",X"52",X"65",X"63",X"6F",X"76",X"65",X"72",X"20",X"73",X"74",X"61",X"73",X"68",
		X"65",X"64",X"20",X"6C",X"6F",X"6F",X"74",X"2E",X"FF",X"63",X"CF",X"00",X"5B",X"6C",X"66",X"5C",
		X"50",X"72",X"6F",X"74",X"65",X"63",X"74",X"20",X"74",X"68",X"65",X"20",X"64",X"72",X"6F",X"70",
		X"70",X"65",X"64",X"5C",X"6C",X"6F",X"6F",X"74",X"2E",X"FF",X"63",X"F0",X"00",X"5E",X"6C",X"66",
		X"5C",X"57",X"61",X"74",X"63",X"68",X"20",X"66",X"6F",X"72",X"20",X"6D",X"75",X"6C",X"74",X"69",
		X"70",X"6C",X"65",X"5C",X"74",X"68",X"65",X"66",X"74",X"73",X"21",X"FF",X"64",X"12",X"00",X"64",
		X"6C",X"66",X"5C",X"54",X"75",X"72",X"6B",X"65",X"79",X"20",X"61",X"69",X"72",X"20",X"72",X"61",
		X"69",X"64",X"21",X"FF",X"64",X"2A",X"00",X"6A",X"6C",X"66",X"5C",X"43",X"79",X"62",X"6F",X"72",
		X"67",X"20",X"74",X"68",X"72",X"65",X"61",X"74",X"21",X"FF",X"64",X"40",X"00",X"67",X"6C",X"66",
		X"5C",X"53",X"68",X"6F",X"70",X"70",X"69",X"6E",X"67",X"20",X"73",X"70",X"72",X"65",X"65",X"21",
		X"FF",X"64",X"57",X"00",X"61",X"6C",X"66",X"5C",X"54",X"75",X"72",X"6B",X"65",X"79",X"73",X"20",
		X"64",X"69",X"73",X"67",X"75",X"69",X"73",X"65",X"64",X"5C",X"61",X"73",X"20",X"62",X"75",X"73",
		X"69",X"6E",X"65",X"73",X"73",X"6D",X"65",X"6E",X"21",X"FF",X"64",X"80",X"00",X"67",X"6C",X"66",
		X"5C",X"4D",X"61",X"6A",X"6F",X"72",X"20",X"61",X"74",X"74",X"61",X"63",X"6B",X"20",X"69",X"73",
		X"5C",X"62",X"72",X"65",X"77",X"69",X"6E",X"67",X"21",X"FF",X"64",X"A0",X"00",X"5E",X"60",X"55",
		X"54",X"75",X"72",X"6B",X"65",X"79",X"73",X"20",X"73",X"75",X"63",X"63",X"65",X"65",X"64",X"2C",
		X"20",X"2D",X"5C",X"5C",X"4E",X"6F",X"20",X"6D",X"6F",X"72",X"65",X"20",X"74",X"72",X"69",X"65",
		X"73",X"2E",X"5C",X"5C",X"47",X"61",X"6D",X"65",X"20",X"6F",X"76",X"65",X"72",X"2E",X"FF",X"64",
		X"D5",X"00",X"5E",X"60",X"55",X"54",X"75",X"72",X"6B",X"65",X"79",X"73",X"20",X"73",X"75",X"63",
		X"63",X"65",X"65",X"64",X"2C",X"20",X"2D",X"5C",X"5C",X"4E",X"6F",X"20",X"6D",X"6F",X"72",X"65",
		X"20",X"74",X"72",X"69",X"65",X"73",X"2E",X"5C",X"5C",X"50",X"6C",X"61",X"79",X"65",X"72",X"20",
		X"31",X"20",X"47",X"61",X"6D",X"65",X"20",X"6F",X"76",X"65",X"72",X"2E",X"FF",X"65",X"13",X"00",
		X"5E",X"60",X"55",X"54",X"75",X"72",X"6B",X"65",X"79",X"73",X"20",X"73",X"75",X"63",X"63",X"65",
		X"65",X"64",X"2C",X"20",X"2D",X"5C",X"5C",X"4E",X"6F",X"20",X"6D",X"6F",X"72",X"65",X"20",X"74",
		X"72",X"69",X"65",X"73",X"2E",X"5C",X"5C",X"50",X"6C",X"61",X"79",X"65",X"72",X"20",X"32",X"20",
		X"47",X"61",X"6D",X"65",X"20",X"6F",X"76",X"65",X"72",X"2E",X"FF",X"65",X"51",X"00",X"58",X"60",
		X"55",X"42",X"6F",X"6E",X"75",X"73",X"20",X"72",X"6F",X"75",X"6E",X"64",X"20",X"65",X"6E",X"64",
		X"65",X"64",X"2C",X"20",X"2D",X"5C",X"5C",X"42",X"79",X"73",X"74",X"61",X"6E",X"64",X"65",X"72",
		X"20",X"64",X"61",X"6D",X"61",X"67",X"65",X"2E",X"FF",X"65",X"7F",X"00",X"55",X"60",X"BB",X"42",
		X"6F",X"6E",X"75",X"73",X"20",X"72",X"6F",X"75",X"6E",X"64",X"20",X"6F",X"76",X"65",X"72",X"2E",
		X"FF",X"65",X"97",X"00",X"76",X"90",X"66",X"35",X"30",X"30",X"30",X"20",X"42",X"4F",X"4E",X"55",
		X"53",X"FF",X"65",X"A8",X"00",X"52",X"60",X"BB",X"43",X"6F",X"6E",X"67",X"72",X"61",X"74",X"75",
		X"6C",X"61",X"74",X"69",X"6F",X"6E",X"73",X"20",X"68",X"65",X"72",X"6F",X"5C",X"6F",X"66",X"20",
		X"68",X"65",X"72",X"6F",X"65",X"73",X"21",X"5C",X"54",X"68",X"65",X"20",X"74",X"75",X"72",X"6B",
		X"65",X"79",X"20",X"74",X"68",X"72",X"65",X"61",X"74",X"20",X"68",X"61",X"73",X"5C",X"65",X"6E",
		X"64",X"65",X"64",X"20",X"66",X"6F",X"72",X"65",X"76",X"65",X"72",X"21",X"5C",X"5C",X"59",X"6F",
		X"75",X"20",X"61",X"72",X"65",X"20",X"72",X"65",X"77",X"61",X"72",X"64",X"65",X"64",X"5C",X"31",
		X"2C",X"30",X"30",X"30",X"2C",X"30",X"30",X"30",X"20",X"62",X"6F",X"6E",X"75",X"73",X"21",X"5C",
		X"54",X"68",X"65",X"20",X"77",X"6F",X"72",X"6C",X"64",X"20",X"69",X"73",X"20",X"66",X"72",X"65",
		X"65",X"2E",X"FF",X"00",X"3A",X"00",X"3A",X"00",X"52",X"00",X"72",X"00",X"92",X"00",X"7A",X"00",
		X"7A",X"00",X"82",X"00",X"C2",X"00",X"A2",X"00",X"8A",X"00",X"72",X"00",X"62",X"00",X"92",X"00",
		X"7A",X"00",X"AA",X"00",X"C2",X"00",X"9A",X"00",X"CA",X"00",X"6A",X"66",X"73",X"66",X"73",X"66",
		X"AD",X"66",X"FF",X"67",X"71",X"68",X"03",X"68",X"7D",X"68",X"F7",X"69",X"79",X"6A",X"3B",X"6A",
		X"DD",X"66",X"FF",X"6B",X"67",X"6B",X"C9",X"68",X"7D",X"6C",X"5B",X"69",X"79",X"6D",X"05",X"6D",
		X"9F",X"6E",X"69",X"00",X"10",X"00",X"20",X"28",X"37",X"8F",X"CC",X"00",X"30",X"FE",X"04",X"00",
		X"00",X"29",X"8C",X"00",X"40",X"FE",X"04",X"00",X"00",X"5D",X"8C",X"00",X"50",X"FE",X"04",X"00",
		X"00",X"2D",X"B4",X"00",X"60",X"FE",X"04",X"00",X"00",X"2D",X"54",X"00",X"70",X"FE",X"04",X"00",
		X"00",X"59",X"9C",X"00",X"80",X"FE",X"04",X"00",X"00",X"35",X"64",X"FF",X"FF",X"00",X"10",X"FE",
		X"20",X"00",X"00",X"00",X"00",X"00",X"20",X"FE",X"20",X"00",X"00",X"00",X"00",X"00",X"30",X"1C",
		X"04",X"01",X"38",X"49",X"9C",X"00",X"40",X"1C",X"04",X"01",X"38",X"49",X"9C",X"00",X"90",X"10",
		X"04",X"34",X"3A",X"49",X"9C",X"00",X"98",X"12",X"04",X"5F",X"3A",X"49",X"9C",X"00",X"A0",X"1C",
		X"06",X"01",X"38",X"49",X"9C",X"00",X"B0",X"1C",X"06",X"01",X"38",X"49",X"9C",X"01",X"10",X"1C",
		X"04",X"01",X"38",X"59",X"5C",X"01",X"30",X"1C",X"04",X"01",X"38",X"51",X"7C",X"FF",X"FF",X"00",
		X"10",X"00",X"02",X"49",X"F8",X"49",X"00",X"00",X"50",X"00",X"02",X"49",X"F8",X"49",X"01",X"00",
		X"90",X"00",X"02",X"49",X"F8",X"49",X"02",X"00",X"D0",X"00",X"02",X"49",X"F8",X"49",X"03",X"01",
		X"10",X"00",X"02",X"49",X"F8",X"49",X"04",X"01",X"30",X"00",X"02",X"49",X"F8",X"49",X"05",X"01",
		X"50",X"00",X"02",X"49",X"F8",X"49",X"06",X"01",X"70",X"00",X"02",X"49",X"F8",X"49",X"07",X"01",
		X"B0",X"00",X"02",X"49",X"F8",X"49",X"08",X"01",X"D0",X"00",X"02",X"49",X"F8",X"49",X"09",X"01",
		X"F0",X"00",X"02",X"49",X"F8",X"49",X"08",X"02",X"10",X"00",X"02",X"49",X"F8",X"49",X"09",X"02",
		X"30",X"00",X"02",X"49",X"F8",X"49",X"08",X"02",X"50",X"00",X"02",X"49",X"F8",X"49",X"09",X"FF",
		X"FF",X"00",X"00",X"14",X"1C",X"01",X"D4",X"48",X"D4",X"00",X"20",X"00",X"20",X"28",X"71",X"48",
		X"CD",X"80",X"50",X"00",X"04",X"48",X"D0",X"38",X"C0",X"80",X"54",X"00",X"04",X"48",X"D0",X"48",
		X"C0",X"80",X"58",X"00",X"04",X"48",X"D0",X"58",X"C0",X"00",X"70",X"FE",X"04",X"00",X"00",X"59",
		X"9C",X"80",X"80",X"1C",X"18",X"01",X"74",X"4D",X"74",X"00",X"90",X"FE",X"06",X"00",X"00",X"35",
		X"64",X"00",X"A0",X"FE",X"06",X"00",X"00",X"4D",X"8C",X"00",X"B0",X"FE",X"04",X"00",X"00",X"75",
		X"BC",X"00",X"E0",X"00",X"04",X"48",X"D0",X"2D",X"54",X"01",X"60",X"FE",X"06",X"00",X"00",X"48",
		X"D0",X"01",X"70",X"FE",X"06",X"00",X"00",X"48",X"D0",X"81",X"80",X"00",X"0A",X"4D",X"71",X"4D",
		X"6C",X"81",X"90",X"00",X"0A",X"4D",X"71",X"4D",X"6C",X"01",X"A0",X"FE",X"06",X"00",X"00",X"48",
		X"D0",X"01",X"B0",X"00",X"36",X"00",X"00",X"AD",X"74",X"02",X"10",X"00",X"38",X"00",X"00",X"F2",
		X"D4",X"FF",X"FF",X"00",X"00",X"16",X"1C",X"8F",X"DC",X"65",X"DC",X"00",X"18",X"00",X"20",X"7E",
		X"B1",X"01",X"39",X"80",X"20",X"1E",X"1A",X"8F",X"64",X"45",X"64",X"00",X"30",X"14",X"0E",X"01",
		X"CC",X"7E",X"B1",X"80",X"50",X"00",X"04",X"65",X"D8",X"55",X"C8",X"80",X"54",X"00",X"04",X"65",
		X"D8",X"65",X"C8",X"80",X"58",X"00",X"04",X"65",X"D8",X"75",X"C8",X"00",X"80",X"16",X"0C",X"8F",
		X"CC",X"59",X"A4",X"00",X"90",X"16",X"0C",X"8F",X"CC",X"49",X"9C",X"81",X"50",X"00",X"04",X"45",
		X"61",X"55",X"51",X"81",X"54",X"00",X"06",X"45",X"5F",X"35",X"51",X"81",X"58",X"00",X"04",X"45",
		X"61",X"45",X"51",X"81",X"5C",X"00",X"06",X"45",X"61",X"4D",X"51",X"01",X"10",X"00",X"3A",X"00",
		X"00",X"F2",X"DC",X"02",X"00",X"00",X"38",X"00",X"00",X"F2",X"64",X"FF",X"FF",X"00",X"10",X"FE",
		X"20",X"00",X"00",X"00",X"00",X"00",X"18",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"FE",
		X"0C",X"00",X"00",X"28",X"80",X"00",X"30",X"FE",X"0C",X"00",X"00",X"60",X"60",X"00",X"40",X"FE",
		X"10",X"00",X"00",X"50",X"60",X"00",X"50",X"FE",X"10",X"00",X"00",X"70",X"80",X"00",X"60",X"FE",
		X"10",X"00",X"00",X"30",X"80",X"00",X"70",X"FE",X"0C",X"00",X"00",X"40",X"A0",X"00",X"80",X"FE",
		X"0C",X"00",X"00",X"58",X"58",X"00",X"90",X"FE",X"10",X"00",X"00",X"78",X"80",X"00",X"A0",X"FE",
		X"0C",X"00",X"00",X"68",X"70",X"80",X"B0",X"16",X"1C",X"8F",X"D4",X"35",X"D4",X"00",X"C0",X"FE",
		X"0C",X"00",X"00",X"30",X"80",X"00",X"D0",X"FE",X"10",X"00",X"00",X"30",X"80",X"00",X"E0",X"FE",
		X"0C",X"00",X"00",X"28",X"80",X"FF",X"FF",X"00",X"10",X"00",X"20",X"6C",X"71",X"01",X"39",X"00",
		X"20",X"00",X"02",X"49",X"F8",X"49",X"00",X"00",X"40",X"FE",X"06",X"00",X"00",X"5D",X"8C",X"00",
		X"50",X"FE",X"04",X"00",X"00",X"29",X"8C",X"00",X"60",X"00",X"02",X"49",X"F8",X"49",X"00",X"00",
		X"70",X"FE",X"04",X"00",X"00",X"2D",X"B4",X"00",X"C0",X"FE",X"04",X"00",X"00",X"2D",X"54",X"00",
		X"E0",X"00",X"02",X"49",X"F8",X"49",X"00",X"01",X"00",X"FE",X"04",X"00",X"00",X"59",X"9C",X"01",
		X"20",X"00",X"02",X"49",X"F8",X"49",X"00",X"01",X"40",X"FE",X"04",X"00",X"00",X"35",X"64",X"01",
		X"90",X"00",X"02",X"49",X"F8",X"49",X"00",X"01",X"E0",X"FE",X"04",X"00",X"00",X"4D",X"8C",X"01",
		X"F0",X"FE",X"04",X"00",X"00",X"75",X"BC",X"02",X"60",X"00",X"02",X"49",X"F8",X"49",X"00",X"02",
		X"E0",X"00",X"02",X"49",X"F8",X"49",X"00",X"FF",X"FF",X"00",X"10",X"00",X"20",X"48",X"38",X"01",
		X"39",X"00",X"20",X"FE",X"06",X"00",X"00",X"3A",X"7A",X"00",X"30",X"FE",X"04",X"00",X"00",X"58",
		X"7A",X"00",X"40",X"00",X"02",X"49",X"F8",X"49",X"00",X"80",X"50",X"1C",X"18",X"01",X"74",X"4D",
		X"74",X"00",X"60",X"FE",X"04",X"00",X"00",X"3A",X"5C",X"00",X"70",X"FE",X"04",X"00",X"00",X"58",
		X"5C",X"00",X"80",X"00",X"02",X"49",X"F8",X"49",X"00",X"00",X"90",X"FE",X"06",X"00",X"00",X"48",
		X"74",X"00",X"A0",X"FE",X"04",X"00",X"00",X"3D",X"64",X"00",X"B0",X"FE",X"04",X"00",X"00",X"51",
		X"6C",X"00",X"C0",X"00",X"02",X"49",X"F8",X"49",X"00",X"00",X"D0",X"00",X"02",X"49",X"F8",X"49",
		X"00",X"00",X"E0",X"FE",X"04",X"00",X"00",X"41",X"64",X"00",X"F0",X"00",X"02",X"49",X"F8",X"49",
		X"00",X"01",X"00",X"FE",X"04",X"00",X"00",X"4D",X"7C",X"81",X"10",X"00",X"0A",X"4D",X"71",X"4D",
		X"38",X"01",X"20",X"00",X"02",X"49",X"F8",X"49",X"00",X"81",X"30",X"00",X"36",X"00",X"00",X"AD",
		X"74",X"01",X"40",X"FE",X"04",X"00",X"00",X"4D",X"5C",X"01",X"50",X"00",X"02",X"49",X"F8",X"49",
		X"00",X"01",X"60",X"FE",X"04",X"00",X"00",X"3A",X"6C",X"01",X"70",X"00",X"02",X"49",X"F8",X"49",
		X"00",X"01",X"80",X"FE",X"04",X"00",X"00",X"55",X"6C",X"FF",X"FF",X"00",X"10",X"FE",X"20",X"00",
		X"00",X"00",X"00",X"00",X"18",X"FE",X"00",X"00",X"00",X"00",X"00",X"80",X"20",X"1C",X"18",X"01",
		X"7C",X"38",X"7C",X"80",X"50",X"1E",X"18",X"8F",X"6C",X"58",X"6C",X"00",X"60",X"14",X"0E",X"01",
		X"CC",X"7E",X"B1",X"00",X"70",X"1E",X"0E",X"8F",X"39",X"6D",X"37",X"81",X"10",X"00",X"0A",X"38",
		X"79",X"13",X"B1",X"81",X"20",X"00",X"0A",X"38",X"79",X"28",X"71",X"81",X"30",X"00",X"0A",X"38",
		X"79",X"16",X"37",X"81",X"40",X"00",X"0A",X"38",X"79",X"28",X"37",X"81",X"50",X"00",X"0A",X"58",
		X"69",X"7E",X"B1",X"81",X"60",X"00",X"0A",X"58",X"69",X"6C",X"71",X"81",X"70",X"00",X"0A",X"58",
		X"69",X"85",X"37",X"81",X"80",X"00",X"0A",X"58",X"69",X"6D",X"37",X"81",X"C0",X"00",X"36",X"00",
		X"00",X"AD",X"7C",X"81",X"D0",X"00",X"36",X"00",X"00",X"F2",X"6C",X"01",X"E0",X"FE",X"06",X"00",
		X"00",X"49",X"7C",X"01",X"F0",X"FE",X"06",X"00",X"00",X"49",X"9C",X"02",X"00",X"FE",X"06",X"00",
		X"00",X"49",X"7C",X"02",X"10",X"FE",X"06",X"00",X"00",X"49",X"9C",X"FF",X"FF",X"00",X"10",X"FE",
		X"20",X"00",X"00",X"00",X"00",X"00",X"18",X"FE",X"20",X"00",X"00",X"00",X"00",X"80",X"20",X"16",
		X"1C",X"8F",X"D0",X"48",X"D0",X"00",X"30",X"FE",X"04",X"00",X"00",X"49",X"7C",X"00",X"40",X"FE",
		X"08",X"00",X"00",X"49",X"7C",X"00",X"50",X"FE",X"04",X"00",X"00",X"49",X"7C",X"00",X"60",X"FE",
		X"06",X"00",X"00",X"49",X"7C",X"80",X"88",X"1E",X"18",X"8F",X"78",X"38",X"78",X"00",X"90",X"FE",
		X"06",X"00",X"00",X"49",X"7C",X"80",X"F0",X"00",X"08",X"48",X"CC",X"48",X"C7",X"81",X"00",X"00",
		X"04",X"48",X"CC",X"48",X"C7",X"81",X"10",X"00",X"04",X"48",X"CC",X"48",X"C7",X"81",X"20",X"00",
		X"3A",X"00",X"00",X"F2",X"D0",X"01",X"30",X"FE",X"06",X"00",X"00",X"49",X"7C",X"01",X"40",X"FE",
		X"06",X"00",X"00",X"49",X"7C",X"81",X"60",X"00",X"0A",X"38",X"75",X"38",X"70",X"81",X"70",X"00",
		X"36",X"00",X"00",X"F2",X"78",X"FF",X"FF",X"00",X"10",X"FE",X"20",X"00",X"00",X"00",X"00",X"00",
		X"20",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"FE",X"08",X"00",X"00",X"28",X"80",X"00",
		X"50",X"FE",X"08",X"00",X"00",X"60",X"60",X"00",X"70",X"FE",X"08",X"00",X"00",X"50",X"60",X"00",
		X"90",X"FE",X"08",X"00",X"00",X"70",X"80",X"00",X"A0",X"FE",X"06",X"00",X"00",X"49",X"7C",X"00",
		X"B0",X"FE",X"08",X"00",X"00",X"30",X"80",X"00",X"C0",X"FE",X"06",X"00",X"00",X"49",X"7C",X"00",
		X"D0",X"FE",X"08",X"00",X"00",X"40",X"A0",X"00",X"E0",X"FE",X"06",X"00",X"00",X"49",X"7C",X"00",
		X"F0",X"FE",X"08",X"00",X"00",X"58",X"58",X"FF",X"FF",X"00",X"10",X"FE",X"20",X"00",X"00",X"00",
		X"00",X"00",X"18",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"16",X"1C",X"8F",X"D4",X"55",
		X"D4",X"00",X"30",X"1C",X"1A",X"01",X"6C",X"65",X"6C",X"80",X"40",X"FE",X"0E",X"00",X"00",X"00",
		X"00",X"80",X"4F",X"FE",X"0E",X"00",X"00",X"00",X"00",X"80",X"5E",X"FE",X"0E",X"00",X"00",X"00",
		X"00",X"80",X"6D",X"FE",X"0E",X"00",X"00",X"00",X"00",X"80",X"7C",X"FE",X"0E",X"00",X"00",X"00",
		X"00",X"80",X"8B",X"FE",X"0E",X"00",X"00",X"00",X"00",X"80",X"E0",X"00",X"04",X"55",X"D0",X"55",
		X"CB",X"80",X"FA",X"FE",X"0E",X"00",X"00",X"00",X"00",X"81",X"00",X"00",X"06",X"65",X"69",X"65",
		X"64",X"81",X"19",X"FE",X"0E",X"00",X"00",X"00",X"00",X"81",X"20",X"00",X"04",X"55",X"D0",X"55",
		X"CB",X"81",X"30",X"00",X"06",X"65",X"69",X"65",X"64",X"81",X"60",X"00",X"38",X"00",X"00",X"AD",
		X"6C",X"81",X"90",X"00",X"3A",X"00",X"00",X"F2",X"6C",X"FF",X"FF",X"00",X"10",X"FE",X"20",X"00",
		X"00",X"00",X"00",X"00",X"30",X"00",X"02",X"49",X"F8",X"49",X"00",X"00",X"50",X"FE",X"04",X"00",
		X"00",X"5D",X"8C",X"00",X"60",X"FE",X"04",X"00",X"00",X"29",X"8C",X"00",X"70",X"00",X"02",X"49",
		X"F8",X"49",X"00",X"00",X"80",X"FE",X"04",X"00",X"00",X"2D",X"B4",X"00",X"D0",X"FE",X"04",X"00",
		X"00",X"2D",X"54",X"00",X"F0",X"00",X"02",X"49",X"F8",X"49",X"00",X"01",X"10",X"FE",X"04",X"00",
		X"00",X"59",X"9C",X"81",X"20",X"1C",X"18",X"01",X"6C",X"35",X"6C",X"01",X"30",X"00",X"02",X"49",
		X"F8",X"49",X"00",X"01",X"50",X"FE",X"04",X"00",X"00",X"35",X"64",X"01",X"80",X"00",X"02",X"49",
		X"F8",X"49",X"00",X"01",X"C0",X"00",X"02",X"49",X"F8",X"49",X"00",X"81",X"D0",X"00",X"0A",X"35",
		X"69",X"35",X"64",X"81",X"E0",X"00",X"0A",X"35",X"69",X"35",X"64",X"01",X"F0",X"FE",X"06",X"00",
		X"00",X"4D",X"8C",X"02",X"00",X"FE",X"04",X"00",X"00",X"75",X"BC",X"02",X"10",X"00",X"36",X"00",
		X"00",X"AD",X"6C",X"02",X"70",X"00",X"02",X"49",X"F8",X"49",X"00",X"02",X"F0",X"00",X"02",X"49",
		X"F8",X"49",X"00",X"FF",X"FF",X"00",X"10",X"FE",X"20",X"00",X"00",X"00",X"00",X"00",X"20",X"FE",
		X"20",X"00",X"00",X"00",X"00",X"00",X"30",X"FE",X"04",X"00",X"00",X"5D",X"8C",X"00",X"40",X"FE",
		X"06",X"00",X"00",X"4D",X"8C",X"00",X"50",X"FE",X"04",X"00",X"00",X"29",X"8C",X"00",X"60",X"FE",
		X"08",X"00",X"00",X"58",X"58",X"00",X"70",X"FE",X"04",X"00",X"00",X"5D",X"8C",X"00",X"80",X"FE",
		X"06",X"00",X"00",X"4D",X"8C",X"00",X"90",X"FE",X"06",X"00",X"00",X"29",X"8C",X"00",X"A0",X"FE",
		X"08",X"00",X"00",X"58",X"58",X"00",X"B0",X"FE",X"06",X"00",X"00",X"5D",X"8C",X"00",X"C0",X"FE",
		X"06",X"00",X"00",X"4D",X"8C",X"00",X"D0",X"FE",X"04",X"00",X"00",X"29",X"8C",X"00",X"E0",X"FE",
		X"08",X"00",X"00",X"58",X"58",X"00",X"F0",X"FE",X"04",X"00",X"00",X"2D",X"B4",X"81",X"30",X"00",
		X"02",X"49",X"F8",X"49",X"00",X"81",X"31",X"00",X"02",X"49",X"F8",X"49",X"00",X"01",X"40",X"FE",
		X"0C",X"00",X"00",X"60",X"60",X"01",X"50",X"FE",X"10",X"00",X"00",X"59",X"9C",X"FF",X"FF",X"00",
		X"10",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"20",X"00",X"00",X"00",X"00",X"00",
		X"12",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"14",X"00",X"30",X"00",X"00",X"00",X"00",X"00",
		X"15",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"16",X"00",X"30",X"00",X"00",X"00",X"00",X"00",
		X"17",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"18",X"00",X"30",X"00",X"00",X"00",X"00",X"00",
		X"19",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"1A",X"00",X"30",X"00",X"00",X"00",X"00",X"00",
		X"1B",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"1C",X"00",X"30",X"00",X"00",X"00",X"00",X"00",
		X"1D",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"1E",X"00",X"30",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"30",X"00",X"00",X"00",X"00",X"00",
		X"21",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"30",X"00",X"00",X"00",X"00",X"00",
		X"23",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"70",X"02",X"04",X"16",X"37",X"00",X"00",X"00",
		X"78",X"04",X"04",X"28",X"37",X"00",X"00",X"00",X"80",X"10",X"04",X"34",X"3A",X"00",X"00",X"00",
		X"88",X"12",X"04",X"5F",X"3A",X"00",X"00",X"00",X"90",X"08",X"04",X"6D",X"37",X"00",X"00",X"00",
		X"98",X"0A",X"04",X"85",X"37",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"2A",X"01",X"44",X"AC",
		X"44",X"00",X"18",X"00",X"20",X"2B",X"44",X"01",X"39",X"00",X"20",X"00",X"20",X"37",X"44",X"01",
		X"CC",X"00",X"28",X"00",X"20",X"43",X"44",X"8F",X"39",X"00",X"30",X"00",X"20",X"4F",X"44",X"8F",
		X"CC",X"00",X"40",X"1C",X"06",X"01",X"38",X"49",X"9C",X"00",X"48",X"1E",X"06",X"8F",X"38",X"49",
		X"9C",X"00",X"50",X"14",X"06",X"01",X"CC",X"49",X"9C",X"80",X"58",X"16",X"06",X"8F",X"CC",X"49",
		X"9C",X"81",X"C0",X"1C",X"06",X"01",X"38",X"49",X"9C",X"01",X"C8",X"1E",X"06",X"8F",X"38",X"49",
		X"9C",X"01",X"D0",X"14",X"06",X"01",X"CC",X"49",X"9C",X"01",X"D8",X"16",X"06",X"8F",X"CC",X"49",
		X"9C",X"FF",X"FF",X"6F",X"0B",X"6F",X"31",X"6F",X"69",X"6F",X"0B",X"6F",X"31",X"6F",X"69",X"6F",
		X"0B",X"6F",X"31",X"6F",X"69",X"6F",X"0B",X"6F",X"31",X"6F",X"69",X"6F",X"0B",X"6F",X"83",X"00",
		X"26",X"00",X"38",X"00",X"1A",X"00",X"26",X"00",X"38",X"00",X"1A",X"00",X"26",X"00",X"38",X"00",
		X"1A",X"00",X"26",X"00",X"38",X"00",X"1A",X"00",X"26",X"00",X"26",X"00",X"2C",X"00",X"00",X"13",
		X"C8",X"00",X"2E",X"00",X"00",X"7A",X"C1",X"00",X"2E",X"00",X"00",X"1A",X"41",X"00",X"30",X"00",
		X"00",X"7A",X"40",X"00",X"30",X"00",X"00",X"05",X"BE",X"00",X"2A",X"48",X"00",X"48",X"1A",X"FF",
		X"FF",X"00",X"2C",X"00",X"00",X"7E",X"C8",X"00",X"2E",X"00",X"00",X"19",X"C1",X"00",X"2E",X"00",
		X"00",X"69",X"41",X"00",X"30",X"00",X"00",X"78",X"C1",X"00",X"30",X"00",X"00",X"18",X"40",X"00",
		X"12",X"FF",X"00",X"3C",X"38",X"00",X"12",X"00",X"00",X"44",X"36",X"00",X"12",X"00",X"00",X"54",
		X"38",X"00",X"2A",X"48",X"00",X"48",X"1A",X"FF",X"FF",X"00",X"2C",X"00",X"00",X"13",X"C8",X"00",
		X"2E",X"00",X"00",X"7A",X"C1",X"00",X"30",X"00",X"00",X"89",X"BF",X"00",X"2A",X"48",X"00",X"48",
		X"1A",X"FF",X"FF",X"00",X"30",X"00",X"00",X"35",X"44",X"00",X"30",X"00",X"00",X"38",X"42",X"00",
		X"12",X"FF",X"00",X"1E",X"3E",X"00",X"12",X"00",X"00",X"26",X"3C",X"00",X"12",X"FF",X"00",X"75",
		X"3E",X"00",X"12",X"00",X"00",X"6A",X"3C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EE",X"60",X"FF",X"FA",X"EE",X"60",X"0F",X"FD",X"F0",X"FE",X"EE",X"60",X"B7",X"8E",X"07",X"5E",
		X"01",X"7E",X"01",X"BD",X"2C",X"50",X"B7",X"6E",X"97",X"BA",X"1E",X"60",X"2F",X"00",X"00",X"00",
		X"0E",X"F0",X"0F",X"F0",X"EE",X"60",X"EC",X"FF",X"EE",X"60",X"ED",X"FE",X"B7",X"8E",X"07",X"5E",
		X"01",X"7E",X"01",X"BD",X"2C",X"50",X"00",X"F0",X"97",X"BA",X"1E",X"60",X"2F",X"00",X"00",X"00",
		X"00",X"00",X"DD",X"F0",X"EE",X"90",X"0F",X"F8",X"0F",X"F8",X"0F",X"F8",X"B7",X"8E",X"07",X"5E",
		X"01",X"7E",X"01",X"BD",X"2C",X"50",X"0F",X"F8",X"97",X"CA",X"1E",X"60",X"2F",X"00",X"00",X"00",
		X"0F",X"FF",X"E0",X"EF",X"EE",X"90",X"FE",X"F0",X"0C",X"EF",X"F3",X"F0",X"B7",X"8E",X"07",X"5E",
		X"01",X"7E",X"01",X"BD",X"2C",X"50",X"00",X"00",X"97",X"BA",X"1E",X"60",X"2F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"B7",X"8E",X"07",X"5E",
		X"01",X"7E",X"01",X"BD",X"2C",X"50",X"00",X"00",X"97",X"BA",X"1E",X"60",X"2F",X"00",X"00",X"00",
		X"00",X"00",X"EE",X"90",X"EE",X"80",X"00",X"00",X"EE",X"90",X"00",X"00",X"B7",X"8E",X"07",X"5E",
		X"01",X"7E",X"01",X"BD",X"2C",X"50",X"00",X"00",X"97",X"BA",X"1E",X"60",X"2F",X"00",X"00",X"00",
		X"00",X"00",X"FE",X"E0",X"EE",X"90",X"AE",X"E9",X"2F",X"51",X"6F",X"C0",X"B7",X"8E",X"07",X"5E",
		X"01",X"7E",X"01",X"BD",X"2C",X"50",X"FF",X"70",X"97",X"BA",X"1E",X"60",X"2F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"B7",X"8E",X"07",X"5E",
		X"01",X"7E",X"01",X"BD",X"2C",X"50",X"00",X"00",X"97",X"BA",X"1E",X"60",X"2F",X"00",X"00",X"00",
		X"EE",X"60",X"FF",X"FA",X"EE",X"60",X"0F",X"FD",X"F0",X"FE",X"EE",X"60",X"B7",X"8E",X"07",X"5E",
		X"01",X"7E",X"01",X"BD",X"2C",X"50",X"B7",X"6E",X"97",X"BA",X"1E",X"60",X"2F",X"00",X"00",X"00",
		X"0E",X"F0",X"0F",X"F0",X"EE",X"60",X"EC",X"FF",X"EE",X"60",X"ED",X"FE",X"B7",X"8E",X"07",X"5E",
		X"01",X"7E",X"01",X"BD",X"2C",X"50",X"00",X"F0",X"97",X"BA",X"1E",X"60",X"2F",X"00",X"00",X"00",
		X"00",X"00",X"DD",X"F0",X"EE",X"90",X"0F",X"F8",X"0F",X"F8",X"0F",X"F8",X"B7",X"8E",X"07",X"5E",
		X"01",X"7E",X"01",X"BD",X"2C",X"50",X"0F",X"F8",X"97",X"CA",X"1E",X"60",X"2F",X"00",X"00",X"00",
		X"0F",X"FF",X"E0",X"EF",X"EE",X"90",X"FE",X"F0",X"0C",X"EF",X"F3",X"F0",X"B7",X"8E",X"07",X"5E",
		X"01",X"7E",X"01",X"BD",X"2C",X"50",X"00",X"00",X"97",X"BA",X"1E",X"60",X"2F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"B7",X"8E",X"07",X"5E",
		X"01",X"7E",X"01",X"BD",X"2C",X"50",X"00",X"00",X"97",X"BA",X"1E",X"60",X"2F",X"00",X"00",X"00",
		X"00",X"00",X"EE",X"40",X"EE",X"80",X"00",X"00",X"EE",X"40",X"00",X"00",X"B7",X"8E",X"07",X"5E",
		X"01",X"7E",X"01",X"BD",X"2C",X"50",X"00",X"00",X"97",X"BA",X"1E",X"60",X"2F",X"00",X"00",X"00",
		X"00",X"00",X"FE",X"E0",X"EE",X"90",X"AE",X"E9",X"2F",X"51",X"6F",X"C0",X"B7",X"8E",X"07",X"5E",
		X"01",X"7E",X"01",X"BD",X"2C",X"50",X"FF",X"70",X"97",X"BA",X"1E",X"60",X"2F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"B7",X"8E",X"07",X"5E",
		X"01",X"7E",X"01",X"BD",X"2C",X"50",X"00",X"00",X"97",X"BA",X"1E",X"60",X"2F",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FA",X"FF",X"0F",X"0F",X"FD",X"F0",X"FE",X"FF",X"0F",X"FF",X"3F",X"DD",X"0D",
		X"FF",X"1F",X"FF",X"4F",X"00",X"00",X"F9",X"FD",X"97",X"8A",X"FF",X"0F",X"22",X"E2",X"00",X"00",
		X"00",X"00",X"0F",X"F0",X"FF",X"0F",X"EC",X"FF",X"FF",X"0F",X"ED",X"FE",X"FF",X"3F",X"DD",X"0D",
		X"FF",X"1F",X"FF",X"4F",X"00",X"00",X"F9",X"FD",X"97",X"8A",X"1E",X"60",X"2F",X"00",X"00",X"00",
		X"00",X"00",X"DD",X"F0",X"FF",X"0F",X"0F",X"F8",X"0F",X"F8",X"0F",X"F8",X"FF",X"3F",X"DD",X"0D",
		X"FF",X"1F",X"FF",X"4F",X"00",X"00",X"0F",X"F8",X"97",X"8A",X"FF",X"0F",X"22",X"E2",X"00",X"00",
		X"00",X"00",X"E0",X"EF",X"FF",X"0F",X"FE",X"F0",X"0C",X"EF",X"F3",X"F0",X"FF",X"3F",X"DD",X"0D",
		X"FF",X"1F",X"FF",X"4F",X"00",X"00",X"00",X"00",X"97",X"8A",X"FF",X"0F",X"22",X"E2",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"3F",X"DD",X"0D",
		X"FF",X"1F",X"FF",X"4F",X"00",X"00",X"00",X"00",X"97",X"8A",X"FF",X"0F",X"22",X"D2",X"00",X"00",
		X"00",X"00",X"FF",X"0F",X"FF",X"0F",X"00",X"00",X"FF",X"0F",X"00",X"00",X"FF",X"3F",X"DD",X"0D",
		X"FF",X"0F",X"FF",X"4F",X"00",X"00",X"00",X"00",X"97",X"8A",X"FF",X"1F",X"22",X"E2",X"00",X"00",
		X"00",X"00",X"FE",X"E1",X"EE",X"90",X"AE",X"E9",X"2F",X"51",X"6F",X"C0",X"FF",X"3F",X"07",X"5E",
		X"01",X"7E",X"01",X"BD",X"01",X"00",X"FF",X"70",X"97",X"BA",X"0F",X"50",X"22",X"E2",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"B7",X"8E",X"07",X"5E",
		X"01",X"7E",X"01",X"BD",X"2C",X"50",X"00",X"00",X"97",X"BA",X"1E",X"60",X"2F",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"BD",X"CA",X"0F",X"F0",X"E0",X"FF",X"BD",X"CA",X"BD",X"40",X"BE",X"1A",
		X"EF",X"1D",X"EF",X"4D",X"2C",X"60",X"0D",X"C8",X"97",X"BA",X"EF",X"3D",X"EF",X"4D",X"00",X"00",
		X"0E",X"F0",X"FC",X"EF",X"BD",X"CA",X"DF",X"EF",X"BD",X"CA",X"CF",X"DF",X"BD",X"40",X"BE",X"1A",
		X"EF",X"1D",X"EF",X"5D",X"2C",X"20",X"0F",X"F0",X"9B",X"B9",X"2F",X"40",X"2F",X"00",X"00",X"00",
		X"00",X"00",X"DD",X"F0",X"EF",X"4F",X"0F",X"F8",X"0F",X"F8",X"0F",X"F8",X"8A",X"60",X"EF",X"4D",
		X"EF",X"0D",X"9D",X"54",X"EF",X"0D",X"0F",X"F8",X"97",X"DA",X"EF",X"3D",X"2F",X"00",X"00",X"00",
		X"0F",X"FF",X"E0",X"EF",X"EF",X"4F",X"FE",X"90",X"0C",X"EF",X"F3",X"F0",X"2C",X"C0",X"EF",X"4D",
		X"EF",X"1D",X"EF",X"3D",X"2C",X"60",X"00",X"00",X"97",X"BA",X"1E",X"60",X"29",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"40",X"EF",X"4F",X"00",X"00",X"00",X"00",X"00",X"00",X"BD",X"40",X"EF",X"4D",
		X"EF",X"6D",X"EF",X"3D",X"7D",X"37",X"00",X"00",X"97",X"BA",X"1E",X"60",X"0F",X"02",X"00",X"00",
		X"00",X"00",X"BD",X"CA",X"BD",X"BA",X"00",X"00",X"BD",X"CA",X"00",X"00",X"BD",X"40",X"EF",X"4D",
		X"EF",X"6D",X"EF",X"3D",X"2C",X"30",X"00",X"00",X"04",X"F0",X"1E",X"40",X"BF",X"20",X"00",X"00",
		X"00",X"00",X"FE",X"E0",X"FE",X"E0",X"AE",X"E9",X"2F",X"51",X"6F",X"C0",X"BD",X"40",X"BD",X"60",
		X"BD",X"80",X"BD",X"90",X"2C",X"50",X"FF",X"70",X"97",X"BA",X"1E",X"60",X"2F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"B7",X"8E",X"07",X"5E",
		X"01",X"7E",X"01",X"BD",X"2C",X"50",X"00",X"00",X"97",X"BA",X"1E",X"60",X"2F",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"CA",X"CD",X"BB",X"0F",X"FD",X"F0",X"EE",X"CD",X"CB",X"FF",X"7F",X"FF",X"0F",
		X"FF",X"4F",X"FF",X"6F",X"2C",X"50",X"B7",X"BE",X"97",X"CA",X"1E",X"60",X"2F",X"00",X"00",X"00",
		X"0E",X"F0",X"0F",X"F0",X"CD",X"AB",X"EC",X"FF",X"CD",X"AB",X"ED",X"FE",X"FF",X"3F",X"FF",X"0F",
		X"FF",X"3F",X"FF",X"5F",X"2C",X"50",X"F9",X"FD",X"97",X"CA",X"1E",X"60",X"2F",X"00",X"00",X"00",
		X"00",X"00",X"DD",X"F0",X"CD",X"AB",X"0F",X"F8",X"0F",X"F8",X"0F",X"F8",X"FF",X"4F",X"FF",X"0F",
		X"FF",X"3F",X"FF",X"5F",X"0E",X"77",X"0F",X"F8",X"97",X"CA",X"1E",X"60",X"2F",X"00",X"00",X"00",
		X"AF",X"FB",X"E0",X"EF",X"CD",X"AB",X"FE",X"F0",X"0C",X"EF",X"F3",X"F0",X"FF",X"7F",X"FF",X"0F",
		X"FF",X"2F",X"FF",X"4F",X"0E",X"67",X"0F",X"EB",X"97",X"BA",X"0A",X"C8",X"0C",X"90",X"00",X"00",
		X"00",X"30",X"F0",X"FF",X"CD",X"AB",X"C0",X"F0",X"0F",X"FF",X"F0",X"F0",X"FF",X"4F",X"FF",X"0F",
		X"FF",X"3F",X"FF",X"5F",X"0E",X"67",X"00",X"10",X"97",X"CA",X"0A",X"C8",X"0C",X"70",X"00",X"00",
		X"00",X"00",X"CD",X"AB",X"CD",X"9B",X"00",X"00",X"CD",X"AB",X"00",X"00",X"FF",X"3F",X"00",X"F0",
		X"FF",X"3F",X"FF",X"5F",X"0F",X"47",X"00",X"00",X"97",X"CA",X"0A",X"C8",X"0C",X"90",X"00",X"00",
		X"00",X"D0",X"FE",X"E0",X"EE",X"90",X"AE",X"E9",X"2F",X"50",X"6F",X"C0",X"FF",X"3F",X"FF",X"0F",
		X"FF",X"3F",X"FF",X"5F",X"2C",X"50",X"FF",X"70",X"97",X"BA",X"1E",X"60",X"2F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"B7",X"8E",X"07",X"5E",
		X"01",X"7E",X"01",X"BD",X"2C",X"50",X"00",X"00",X"97",X"BA",X"1E",X"60",X"2F",X"00",X"00",X"00",
		X"45",X"06",X"DF",X"90",X"75",X"12",X"AA",X"AA",X"AA",X"25",X"29",X"28",X"78",X"45",X"45",X"45",
		X"45",X"07",X"5F",X"10",X"79",X"11",X"2A",X"2A",X"2A",X"24",X"23",X"22",X"76",X"45",X"45",X"45",
		X"45",X"49",X"08",X"47",X"71",X"7A",X"46",X"7C",X"7D",X"72",X"27",X"26",X"77",X"45",X"45",X"45",
		X"45",X"C9",X"09",X"C7",X"59",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
		X"45",X"5D",X"43",X"42",X"58",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
		X"45",X"45",X"04",X"41",X"5B",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
		X"45",X"45",X"05",X"C1",X"DB",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
		X"45",X"45",X"C3",X"C2",X"D8",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
		X"45",X"0C",X"44",X"4A",X"D9",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
		X"45",X"CD",X"C4",X"CA",X"F1",X"FA",X"C6",X"9A",X"FD",X"F2",X"A7",X"A6",X"F7",X"45",X"45",X"45",
		X"45",X"4E",X"0D",X"54",X"F9",X"AA",X"19",X"16",X"AA",X"A4",X"A3",X"A2",X"F8",X"45",X"45",X"45",
		X"45",X"CE",X"0E",X"D4",X"F5",X"2A",X"18",X"17",X"2A",X"A5",X"9E",X"9D",X"F8",X"45",X"45",X"45",
		X"45",X"C9",X"C4",X"10",X"35",X"45",X"45",X"45",X"74",X"25",X"29",X"28",X"78",X"45",X"45",X"45",
		X"45",X"BA",X"B8",X"BB",X"B5",X"45",X"45",X"45",X"74",X"24",X"23",X"22",X"78",X"45",X"45",X"45",
		X"45",X"45",X"B9",X"B7",X"B4",X"45",X"45",X"73",X"7D",X"72",X"27",X"26",X"77",X"45",X"45",X"45",
		X"45",X"45",X"B6",X"F0",X"EF",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
		X"45",X"67",X"69",X"68",X"6B",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
		X"45",X"65",X"64",X"63",X"6A",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
		X"45",X"E5",X"E4",X"E3",X"EA",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
		X"45",X"E7",X"E9",X"66",X"6C",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
		X"45",X"45",X"36",X"70",X"6F",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
		X"45",X"45",X"39",X"37",X"34",X"45",X"45",X"F3",X"FD",X"F2",X"A7",X"A6",X"F7",X"45",X"45",X"45",
		X"45",X"3A",X"38",X"3B",X"35",X"45",X"45",X"45",X"F4",X"A4",X"A3",X"A2",X"F8",X"45",X"45",X"45",
		X"45",X"C9",X"08",X"47",X"B5",X"45",X"45",X"45",X"F4",X"A5",X"9E",X"9D",X"78",X"45",X"45",X"45",
		X"45",X"02",X"AB",X"81",X"5B",X"45",X"D7",X"7B",X"BE",X"25",X"29",X"28",X"78",X"45",X"45",X"45",
		X"45",X"20",X"2B",X"01",X"5B",X"45",X"D7",X"7E",X"3E",X"24",X"23",X"22",X"76",X"45",X"45",X"45",
		X"45",X"45",X"3D",X"2C",X"5B",X"45",X"53",X"48",X"7D",X"72",X"27",X"26",X"77",X"45",X"45",X"45",
		X"45",X"45",X"3C",X"AC",X"59",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
		X"45",X"45",X"43",X"42",X"58",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
		X"45",X"45",X"04",X"41",X"5B",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
		X"45",X"45",X"05",X"C1",X"DB",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
		X"45",X"CD",X"C3",X"C2",X"D8",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
		X"45",X"6D",X"13",X"15",X"D9",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
		X"45",X"0B",X"93",X"95",X"5B",X"45",X"D3",X"C8",X"FD",X"F2",X"A7",X"A6",X"F7",X"45",X"45",X"45",
		X"45",X"40",X"5A",X"5C",X"5B",X"45",X"57",X"0A",X"BE",X"A4",X"A3",X"A2",X"F8",X"45",X"45",X"45",
		X"45",X"C0",X"3F",X"DC",X"5B",X"45",X"57",X"51",X"3E",X"A5",X"9E",X"9D",X"F8",X"45",X"45",X"45",
		X"45",X"45",X"44",X"90",X"75",X"55",X"83",X"83",X"83",X"25",X"29",X"28",X"78",X"45",X"45",X"45",
		X"45",X"0F",X"C4",X"10",X"79",X"56",X"03",X"03",X"03",X"24",X"23",X"22",X"78",X"45",X"45",X"45",
		X"45",X"45",X"1C",X"94",X"71",X"7A",X"46",X"48",X"7D",X"72",X"27",X"26",X"77",X"45",X"45",X"45",
		X"45",X"45",X"1F",X"14",X"59",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
		X"45",X"45",X"2F",X"21",X"58",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
		X"45",X"45",X"2E",X"2D",X"5B",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
		X"45",X"45",X"AE",X"AD",X"5B",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
		X"45",X"45",X"AF",X"A1",X"D8",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
		X"45",X"4C",X"44",X"30",X"D9",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
		X"45",X"52",X"C4",X"B0",X"F1",X"FA",X"C6",X"C8",X"FD",X"F2",X"A7",X"A6",X"F7",X"45",X"45",X"45",
		X"45",X"5E",X"60",X"54",X"F9",X"83",X"1B",X"4B",X"83",X"A4",X"A3",X"A2",X"F6",X"45",X"45",X"45",
		X"45",X"DE",X"C4",X"D4",X"F5",X"03",X"03",X"03",X"03",X"A5",X"9E",X"9D",X"F8",X"45",X"45",X"45",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"21",X"21",X"1D",
		X"1D",X"1D",X"1D",X"1C",X"1C",X"1C",X"1C",X"1C",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1A",X"1A",
		X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"21",X"21",X"1D",
		X"1D",X"1D",X"1D",X"1C",X"1C",X"1C",X"1C",X"1C",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1A",X"1A",
		X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"21",X"21",X"1D",
		X"1D",X"1D",X"1D",X"1C",X"1C",X"1C",X"1C",X"1C",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1A",X"1A",
		X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"21",X"21",X"1D",
		X"1D",X"1D",X"1D",X"1C",X"1C",X"1C",X"1C",X"1C",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1A",X"1A",
		X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"72",
		X"72",X"72",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"70",X"70",X"70",X"70",X"70",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"71",X"71",X"75",
		X"75",X"75",X"75",X"76",X"76",X"76",X"76",X"76",X"77",X"77",X"77",X"77",X"77",X"77",X"78",X"78",
		X"78",X"78",X"78",X"78",X"78",X"78",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"70",X"70",X"70",X"70",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"71",X"71",X"75",
		X"75",X"75",X"75",X"76",X"76",X"76",X"76",X"76",X"77",X"77",X"77",X"77",X"77",X"77",X"78",X"78",
		X"78",X"78",X"78",X"78",X"78",X"78",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",
		X"8A",X"8A",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"88",X"88",X"88",X"88",X"88",
		X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"71",X"71",X"75",
		X"75",X"75",X"75",X"76",X"76",X"76",X"76",X"76",X"77",X"77",X"77",X"77",X"77",X"77",X"78",X"78",
		X"78",X"78",X"78",X"78",X"78",X"78",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",
		X"8A",X"8A",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"88",X"88",X"88",X"88",X"88",
		X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"71",X"71",X"75",
		X"75",X"75",X"75",X"76",X"76",X"76",X"76",X"76",X"77",X"77",X"77",X"77",X"77",X"77",X"78",X"78",
		X"78",X"78",X"78",X"78",X"78",X"78",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
