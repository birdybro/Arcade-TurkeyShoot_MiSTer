library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity turkey_shoot_graph2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of turkey_shoot_graph2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"FF",
		X"AF",X"F2",X"22",X"FF",X"2A",X"22",X"CC",X"2F",X"EE",X"DD",X"EA",X"EE",X"E2",X"EE",X"EE",X"2C",
		X"C2",X"77",X"CC",X"22",X"AA",X"CC",X"EE",X"AA",X"AA",X"CC",X"AA",X"AA",X"7F",X"CC",X"77",X"FA",
		X"CC",X"CC",X"CC",X"CC",X"88",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"66",X"66",X"66",X"66",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"3F",X"FF",X"FF",X"F3",X"FF",X"FF",X"F3",X"F3",X"FF",X"FF",X"F3",X"33",X"FF",
		X"FF",X"F3",X"F3",X"FF",X"FF",X"FF",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"FF",X"FF",X"FF",X"FF",
		X"77",X"77",X"77",X"F7",X"77",X"77",X"77",X"F7",X"77",X"77",X"77",X"F7",X"77",X"77",X"77",X"F7",
		X"77",X"77",X"77",X"F7",X"77",X"77",X"77",X"F7",X"77",X"77",X"77",X"F7",X"77",X"77",X"77",X"F7",
		X"77",X"77",X"77",X"F7",X"77",X"77",X"77",X"F7",X"77",X"77",X"77",X"F7",X"77",X"77",X"77",X"F7",
		X"77",X"77",X"77",X"F7",X"77",X"77",X"77",X"F7",X"FF",X"FF",X"FF",X"FF",X"77",X"77",X"77",X"F7",
		X"77",X"FF",X"7F",X"CF",X"99",X"FF",X"9C",X"9C",X"88",X"FC",X"88",X"88",X"77",X"57",X"55",X"75",
		X"77",X"57",X"75",X"5C",X"57",X"57",X"75",X"5C",X"75",X"77",X"75",X"75",X"88",X"88",X"88",X"88",
		X"99",X"99",X"99",X"99",X"88",X"88",X"88",X"88",X"77",X"77",X"77",X"7C",X"77",X"77",X"77",X"7C",
		X"77",X"77",X"77",X"72",X"8A",X"8A",X"8A",X"A2",X"8A",X"8A",X"8A",X"A2",X"8A",X"8A",X"8A",X"A2",
		X"77",X"77",X"77",X"FF",X"99",X"F9",X"99",X"F9",X"88",X"88",X"88",X"88",X"57",X"75",X"75",X"77",
		X"27",X"75",X"7F",X"77",X"27",X"55",X"75",X"77",X"57",X"75",X"75",X"55",X"88",X"88",X"FF",X"88",
		X"F9",X"99",X"CF",X"99",X"88",X"88",X"8C",X"88",X"C7",X"77",X"77",X"77",X"C7",X"77",X"77",X"77",
		X"27",X"77",X"77",X"77",X"2A",X"A8",X"A8",X"A8",X"2A",X"A8",X"A8",X"A8",X"2A",X"A8",X"A8",X"A8",
		X"FF",X"FF",X"FF",X"FF",X"DD",X"FF",X"FF",X"DD",X"FD",X"DF",X"DF",X"DD",X"FF",X"DD",X"DD",X"DD",
		X"DD",X"FD",X"F3",X"DD",X"ED",X"33",X"3F",X"33",X"ED",X"FF",X"FF",X"FF",X"DE",X"F1",X"F1",X"F1",
		X"DD",X"F1",X"F1",X"1F",X"DD",X"F1",X"F1",X"1F",X"EE",X"F1",X"F1",X"1F",X"DD",X"F1",X"F1",X"1F",
		X"ED",X"F1",X"F1",X"1F",X"DF",X"F1",X"FF",X"F1",X"DD",X"FF",X"F3",X"FF",X"FD",X"33",X"3E",X"33",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"DF",X"FF",X"FF",
		X"33",X"DD",X"33",X"FF",X"FF",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"1F",X"FF",
		X"FF",X"F1",X"FF",X"FF",X"FF",X"F1",X"FF",X"FF",X"11",X"F1",X"1F",X"EF",X"FF",X"F1",X"1F",X"EE",
		X"FF",X"F1",X"FF",X"ED",X"FF",X"1F",X"FF",X"DD",X"33",X"FF",X"33",X"DD",X"DD",X"33",X"EE",X"DD",
		X"77",X"77",X"77",X"1B",X"B1",X"B1",X"B1",X"22",X"22",X"22",X"22",X"22",X"21",X"11",X"11",X"12",
		X"12",X"F1",X"FF",X"F1",X"21",X"21",X"11",X"12",X"2F",X"21",X"FF",X"F1",X"11",X"21",X"F2",X"21",
		X"2F",X"22",X"F2",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"B1",X"B1",X"B1",X"B1",
		X"77",X"FF",X"FF",X"77",X"77",X"AA",X"AA",X"77",X"99",X"AC",X"AC",X"99",X"99",X"AC",X"AC",X"99",
		X"B1",X"77",X"77",X"88",X"22",X"B1",X"B1",X"B1",X"22",X"22",X"22",X"22",X"11",X"11",X"11",X"22",
		X"FF",X"1F",X"FF",X"12",X"11",X"1F",X"11",X"F2",X"F2",X"1F",X"FF",X"22",X"F2",X"11",X"11",X"12",
		X"F2",X"2F",X"FF",X"2F",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"B1",X"B1",X"B1",X"B1",
		X"77",X"FF",X"FF",X"77",X"77",X"AA",X"AA",X"79",X"99",X"CA",X"CA",X"99",X"99",X"CA",X"CA",X"99",
		X"66",X"22",X"22",X"F7",X"FF",X"2C",X"22",X"F7",X"77",X"2C",X"0C",X"F0",X"77",X"2C",X"0C",X"07",
		X"77",X"2C",X"C2",X"07",X"77",X"2C",X"22",X"00",X"77",X"2C",X"CC",X"07",X"66",X"00",X"00",X"F7",
		X"66",X"78",X"77",X"77",X"FF",X"22",X"4C",X"F7",X"77",X"22",X"4C",X"47",X"77",X"22",X"C2",X"47",
		X"77",X"22",X"22",X"47",X"77",X"CC",X"CC",X"47",X"77",X"44",X"44",X"F7",X"66",X"CC",X"CC",X"F7",
		X"FF",X"1F",X"77",X"7F",X"FF",X"F1",X"07",X"7F",X"FF",X"F1",X"07",X"7F",X"FF",X"F1",X"07",X"78",
		X"FF",X"F1",X"07",X"78",X"11",X"17",X"07",X"78",X"FF",X"F7",X"07",X"78",X"F4",X"44",X"07",X"78",
		X"F4",X"F7",X"07",X"78",X"F4",X"47",X"07",X"78",X"F4",X"77",X"07",X"78",X"74",X"44",X"07",X"78",
		X"07",X"77",X"07",X"78",X"07",X"77",X"07",X"78",X"0D",X"77",X"07",X"DE",X"F9",X"22",X"F2",X"96",
		X"F0",X"00",X"FF",X"FF",X"0F",X"FF",X"FF",X"FF",X"FF",X"1F",X"FF",X"FF",X"F1",X"F1",X"FF",X"FF",
		X"F1",X"FF",X"FF",X"FF",X"FF",X"1F",X"FF",X"FF",X"FF",X"F1",X"FF",X"FF",X"FF",X"F1",X"FF",X"FF",
		X"F1",X"F1",X"FF",X"FF",X"FF",X"1F",X"FF",X"FF",X"0F",X"FF",X"FF",X"FF",X"F0",X"F0",X"FF",X"FF",
		X"FF",X"0F",X"FF",X"FF",X"F9",X"77",X"FF",X"FF",X"F9",X"77",X"FF",X"FF",X"FF",X"8F",X"FF",X"FF",
		X"99",X"AA",X"AA",X"AA",X"99",X"CC",X"CC",X"AC",X"99",X"CC",X"2C",X"AC",X"99",X"C2",X"3C",X"32",
		X"99",X"22",X"33",X"32",X"99",X"C2",X"32",X"32",X"99",X"C2",X"3C",X"32",X"99",X"C2",X"3C",X"32",
		X"99",X"CC",X"3C",X"32",X"99",X"CC",X"CC",X"AC",X"88",X"88",X"88",X"88",X"EE",X"EE",X"0E",X"E0",
		X"EE",X"EE",X"0E",X"E0",X"EE",X"EE",X"0E",X"EE",X"88",X"88",X"88",X"88",X"77",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"99",X"CA",X"CC",X"CC",X"99",X"CA",X"CC",X"2C",X"99",X"23",X"C3",X"2C",X"99",
		X"23",X"32",X"22",X"99",X"23",X"23",X"22",X"99",X"23",X"C2",X"2C",X"99",X"23",X"C2",X"2C",X"99",
		X"23",X"33",X"CC",X"99",X"CA",X"CC",X"CC",X"99",X"00",X"08",X"E8",X"88",X"EE",X"E0",X"EE",X"EE",
		X"00",X"E0",X"EE",X"EE",X"EE",X"0E",X"0E",X"EE",X"88",X"88",X"88",X"88",X"AA",X"AA",X"AA",X"AA",
		X"F9",X"FF",X"FF",X"9F",X"F9",X"FF",X"FF",X"91",X"F9",X"77",X"77",X"17",X"F9",X"77",X"71",X"91",
		X"F1",X"71",X"71",X"97",X"F1",X"71",X"77",X"97",X"F1",X"71",X"77",X"77",X"F1",X"91",X"99",X"99",
		X"F1",X"77",X"73",X"77",X"FF",X"99",X"99",X"99",X"FF",X"77",X"77",X"77",X"99",X"99",X"99",X"99",
		X"F7",X"37",X"37",X"37",X"99",X"93",X"39",X"99",X"F7",X"73",X"37",X"77",X"F7",X"37",X"77",X"77",
		X"CC",X"CC",X"CA",X"AA",X"CC",X"CC",X"CA",X"CA",X"4C",X"44",X"4A",X"4A",X"4C",X"44",X"4A",X"4E",
		X"4C",X"44",X"4A",X"4E",X"4C",X"44",X"4A",X"4E",X"4C",X"44",X"4A",X"4E",X"4C",X"4C",X"4A",X"AE",
		X"CC",X"CC",X"CA",X"4E",X"CC",X"CC",X"9A",X"4E",X"99",X"99",X"8A",X"4E",X"77",X"77",X"8A",X"CE",
		X"77",X"77",X"8A",X"CE",X"77",X"77",X"8A",X"DE",X"88",X"88",X"CC",X"CC",X"66",X"66",X"66",X"66",
		X"88",X"88",X"88",X"8C",X"F7",X"33",X"7B",X"CF",X"FF",X"E3",X"BB",X"CC",X"3F",X"3F",X"BB",X"B7",
		X"3F",X"3F",X"BB",X"B7",X"33",X"F2",X"BB",X"BB",X"33",X"C2",X"BB",X"BF",X"33",X"2F",X"BB",X"99",
		X"33",X"FB",X"FB",X"FF",X"73",X"BB",X"CF",X"CC",X"73",X"FB",X"22",X"C7",X"73",X"2B",X"FF",X"F7",
		X"73",X"2F",X"BB",X"F7",X"73",X"CF",X"BB",X"F7",X"73",X"F2",X"BB",X"F7",X"73",X"22",X"FF",X"F7",
		X"88",X"88",X"88",X"88",X"55",X"55",X"44",X"77",X"55",X"55",X"44",X"CC",X"55",X"55",X"4F",X"FF",
		X"FF",X"FF",X"F2",X"4F",X"F7",X"CC",X"22",X"44",X"F7",X"C2",X"C2",X"44",X"F7",X"22",X"22",X"44",
		X"F7",X"22",X"F2",X"F4",X"F7",X"22",X"4F",X"7F",X"F7",X"22",X"44",X"7F",X"F7",X"22",X"44",X"74",
		X"F7",X"CC",X"44",X"44",X"F7",X"C2",X"24",X"44",X"F7",X"F2",X"22",X"4F",X"F7",X"22",X"22",X"77",
		X"ED",X"CF",X"CC",X"DF",X"77",X"CF",X"CC",X"7F",X"77",X"CF",X"CC",X"7F",X"87",X"CF",X"CC",X"7F",
		X"89",X"CF",X"CC",X"9F",X"89",X"CF",X"C2",X"9F",X"89",X"CF",X"22",X"9F",X"89",X"2F",X"22",X"9F",
		X"89",X"2F",X"22",X"9F",X"ED",X"2F",X"22",X"DF",X"89",X"2F",X"22",X"9F",X"89",X"2F",X"22",X"9F",
		X"89",X"2F",X"22",X"9F",X"89",X"2F",X"22",X"9F",X"ED",X"2F",X"22",X"DF",X"69",X"2F",X"22",X"9F",
		X"CC",X"AA",X"CA",X"CC",X"CC",X"AC",X"CA",X"CC",X"22",X"A2",X"2A",X"22",X"22",X"A2",X"2A",X"22",
		X"22",X"A2",X"2A",X"22",X"22",X"A2",X"2A",X"22",X"22",X"A2",X"2A",X"22",X"2C",X"AA",X"2A",X"22",
		X"CC",X"A2",X"CA",X"CC",X"CC",X"A2",X"CA",X"99",X"99",X"A2",X"F9",X"98",X"77",X"A2",X"F7",X"78",
		X"77",X"A2",X"F7",X"78",X"77",X"AA",X"F7",X"78",X"88",X"CC",X"C8",X"8C",X"66",X"66",X"66",X"66",
		X"89",X"2F",X"22",X"97",X"89",X"2F",X"22",X"97",X"89",X"2F",X"22",X"97",X"89",X"2F",X"22",X"97",
		X"89",X"2F",X"22",X"97",X"89",X"2F",X"22",X"97",X"89",X"2F",X"22",X"97",X"89",X"F2",X"FF",X"97",
		X"89",X"FF",X"FF",X"97",X"ED",X"2F",X"22",X"D7",X"89",X"AE",X"AA",X"97",X"89",X"F7",X"77",X"97",
		X"89",X"F7",X"77",X"97",X"89",X"F7",X"77",X"9C",X"89",X"77",X"CC",X"97",X"66",X"66",X"66",X"66",
		X"9F",X"12",X"21",X"F7",X"FF",X"11",X"21",X"F7",X"11",X"21",X"12",X"11",X"77",X"22",X"2C",X"F7",
		X"79",X"4C",X"CC",X"F9",X"7F",X"EE",X"EE",X"FF",X"7F",X"98",X"77",X"94",X"7F",X"74",X"77",X"77",
		X"7F",X"42",X"22",X"F7",X"77",X"42",X"24",X"F7",X"77",X"42",X"24",X"F7",X"77",X"44",X"24",X"F7",
		X"44",X"E4",X"42",X"44",X"FF",X"E2",X"22",X"F7",X"7F",X"22",X"22",X"F7",X"7F",X"22",X"22",X"F7",
		X"1F",X"12",X"22",X"F9",X"1F",X"12",X"22",X"FF",X"11",X"22",X"22",X"77",X"7F",X"C2",X"22",X"77",
		X"4F",X"CC",X"C2",X"97",X"F4",X"EE",X"EE",X"F7",X"99",X"47",X"79",X"F7",X"77",X"47",X"77",X"F7",
		X"4F",X"22",X"22",X"F7",X"4F",X"22",X"22",X"77",X"4F",X"42",X"22",X"77",X"4F",X"42",X"22",X"77",
		X"44",X"22",X"2E",X"99",X"7F",X"22",X"2E",X"FF",X"7F",X"22",X"22",X"F7",X"7F",X"22",X"22",X"F7",
		X"0F",X"22",X"22",X"F9",X"70",X"22",X"22",X"FF",X"7F",X"02",X"22",X"77",X"7F",X"02",X"22",X"77",
		X"0F",X"CC",X"C2",X"97",X"0F",X"EE",X"EE",X"F7",X"09",X"07",X"79",X"F7",X"07",X"07",X"77",X"F7",
		X"00",X"22",X"22",X"F7",X"7F",X"22",X"22",X"77",X"1F",X"22",X"22",X"77",X"71",X"22",X"22",X"77",
		X"7F",X"12",X"2E",X"99",X"7F",X"12",X"2E",X"FF",X"1F",X"22",X"22",X"F7",X"1F",X"22",X"22",X"F7",
		X"9F",X"02",X"22",X"F7",X"FF",X"22",X"22",X"F7",X"77",X"22",X"22",X"F0",X"77",X"20",X"22",X"F7",
		X"79",X"0C",X"C2",X"F7",X"7F",X"0E",X"E0",X"F7",X"7F",X"07",X"70",X"97",X"7F",X"00",X"70",X"77",
		X"00",X"20",X"02",X"00",X"77",X"22",X"22",X"F7",X"77",X"12",X"22",X"F7",X"77",X"22",X"22",X"F7",
		X"99",X"E2",X"22",X"F1",X"FF",X"E1",X"22",X"F7",X"7F",X"12",X"22",X"F7",X"7F",X"12",X"21",X"F7",
		X"8A",X"77",X"8F",X"FF",X"AA",X"77",X"8F",X"FF",X"FE",X"F6",X"66",X"66",X"FA",X"77",X"77",X"77",
		X"FA",X"33",X"37",X"33",X"FC",X"77",X"37",X"73",X"FF",X"73",X"37",X"38",X"F8",X"73",X"37",X"33",
		X"C8",X"77",X"77",X"77",X"7F",X"33",X"33",X"33",X"7F",X"98",X"8F",X"FF",X"7F",X"98",X"8F",X"FF",
		X"7F",X"EA",X"8F",X"FF",X"7F",X"DC",X"EA",X"FF",X"7F",X"DE",X"DA",X"FF",X"7F",X"DD",X"DA",X"FF",
		X"7F",X"73",X"77",X"77",X"7F",X"73",X"77",X"77",X"74",X"73",X"77",X"77",X"74",X"7F",X"77",X"77",
		X"74",X"73",X"77",X"77",X"4F",X"73",X"77",X"77",X"4F",X"73",X"77",X"77",X"7F",X"7F",X"77",X"77",
		X"7F",X"73",X"77",X"77",X"7F",X"73",X"77",X"77",X"7F",X"73",X"77",X"77",X"4F",X"7F",X"77",X"77",
		X"4F",X"73",X"77",X"77",X"44",X"7F",X"77",X"77",X"44",X"FF",X"FF",X"FF",X"7F",X"70",X"77",X"77",
		X"8C",X"FF",X"FF",X"FB",X"77",X"FF",X"11",X"FF",X"77",X"CC",X"1F",X"F1",X"77",X"77",X"1F",X"F1",
		X"77",X"99",X"19",X"F1",X"77",X"88",X"18",X"71",X"77",X"88",X"18",X"71",X"77",X"88",X"1F",X"91",
		X"7F",X"88",X"18",X"81",X"7F",X"88",X"18",X"F1",X"7F",X"88",X"18",X"81",X"FF",X"FF",X"FF",X"FF",
		X"B8",X"88",X"8B",X"B8",X"B9",X"99",X"9B",X"B9",X"B8",X"88",X"8B",X"B8",X"FF",X"FF",X"FF",X"FF",
		X"11",X"11",X"11",X"7F",X"11",X"11",X"11",X"7F",X"11",X"C1",X"11",X"7F",X"C1",X"1C",X"C1",X"7F",
		X"1C",X"11",X"11",X"7F",X"CC",X"CF",X"CC",X"7F",X"99",X"F9",X"99",X"7F",X"88",X"F8",X"88",X"7F",
		X"88",X"FF",X"88",X"7F",X"88",X"CC",X"88",X"7F",X"88",X"88",X"88",X"7F",X"FF",X"FF",X"FF",X"7F",
		X"66",X"76",X"66",X"66",X"66",X"66",X"66",X"66",X"E6",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"FF",X"FF",X"FF",X"FF",X"77",X"77",X"77",X"7F",X"CC",X"CC",X"CC",X"7F",X"CC",X"CC",X"CC",X"7F",
		X"CC",X"CC",X"CC",X"7F",X"CC",X"CC",X"CC",X"7F",X"11",X"11",X"11",X"7F",X"11",X"11",X"11",X"7F",
		X"11",X"11",X"11",X"7F",X"11",X"11",X"11",X"7F",X"11",X"1C",X"11",X"7F",X"1C",X"11",X"11",X"7F",
		X"11",X"11",X"C1",X"7F",X"11",X"11",X"1C",X"7F",X"C1",X"11",X"11",X"7F",X"1C",X"11",X"C1",X"7F",
		X"BF",X"FF",X"FF",X"FF",X"FB",X"FF",X"FF",X"FF",X"FF",X"BB",X"FF",X"FF",X"F1",X"FF",X"BF",X"FF",
		X"1F",X"11",X"7B",X"FF",X"1F",X"88",X"77",X"FF",X"19",X"88",X"17",X"FF",X"18",X"88",X"17",X"11",
		X"18",X"88",X"17",X"17",X"18",X"88",X"77",X"77",X"81",X"11",X"17",X"11",X"FF",X"FF",X"FF",X"FF",
		X"B8",X"8B",X"B8",X"8B",X"B9",X"9B",X"B9",X"9B",X"B8",X"8B",X"B8",X"8B",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"33",X"FF",X"FF",X"FF",X"F3",X"F3",X"3F",X"FF",X"F3",X"3F",X"FF",X"FF",X"F3",X"F3",X"3F",X"FF",
		X"F3",X"FF",X"FF",X"FF",X"FF",X"33",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"F1",X"FF",X"FF",
		X"F1",X"1F",X"FF",X"FF",X"F1",X"F1",X"FF",X"FF",X"F1",X"FF",X"FF",X"FF",X"F1",X"11",X"FF",X"FF",
		X"77",X"FA",X"AF",X"FE",X"7C",X"FA",X"AC",X"FE",X"7C",X"FA",X"CF",X"FC",X"72",X"FF",X"FC",X"CF",
		X"72",X"FF",X"CF",X"FC",X"72",X"FF",X"CF",X"CF",X"72",X"FF",X"FC",X"FC",X"72",X"FF",X"FC",X"CF",
		X"77",X"AA",X"9F",X"EC",X"77",X"AE",X"AC",X"CF",X"77",X"CF",X"AA",X"AA",X"77",X"FF",X"AA",X"AA",
		X"7C",X"FF",X"AA",X"AA",X"6C",X"FF",X"AA",X"AA",X"FF",X"F6",X"E2",X"2E",X"FF",X"66",X"66",X"66",
		X"9F",X"A7",X"C2",X"88",X"9F",X"A7",X"22",X"88",X"9F",X"A7",X"22",X"88",X"9F",X"E7",X"22",X"88",
		X"9F",X"E7",X"22",X"88",X"9F",X"E7",X"77",X"F8",X"FF",X"E7",X"87",X"C8",X"CF",X"D7",X"77",X"88",
		X"9F",X"E6",X"66",X"88",X"9F",X"66",X"66",X"88",X"9F",X"66",X"66",X"88",X"FF",X"66",X"66",X"FF",
		X"66",X"66",X"66",X"66",X"66",X"A6",X"88",X"67",X"66",X"AA",X"66",X"66",X"66",X"6A",X"66",X"66",
		X"7F",X"77",X"88",X"88",X"7F",X"88",X"99",X"88",X"7F",X"AF",X"CC",X"F8",X"7F",X"A7",X"CC",X"88",
		X"7F",X"A7",X"CC",X"88",X"7F",X"A7",X"CC",X"88",X"7F",X"A7",X"CC",X"88",X"FF",X"A7",X"CC",X"F8",
		X"8F",X"A7",X"CC",X"C8",X"9F",X"A7",X"C7",X"88",X"9F",X"A7",X"ED",X"88",X"FF",X"A7",X"C7",X"88",
		X"CF",X"A7",X"C7",X"88",X"9F",X"A7",X"C7",X"88",X"9F",X"A7",X"CC",X"F8",X"9F",X"A7",X"CC",X"88",
		X"7F",X"7F",X"7F",X"F7",X"7F",X"7F",X"7F",X"F7",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"77",X"77",X"77",X"77",X"EE",X"EE",X"EE",X"E7",X"EE",X"EE",X"EE",X"E7",X"EE",X"EE",X"EE",X"DD",
		X"EE",X"EE",X"EE",X"E7",X"EE",X"EE",X"EE",X"DD",X"EE",X"EE",X"EE",X"E7",X"EE",X"EE",X"EE",X"DD",
		X"EE",X"EE",X"EE",X"E7",X"EE",X"EE",X"EE",X"E7",X"77",X"77",X"77",X"77",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"7F",X"F7",X"F7",X"7F",X"7F",X"F7",X"F7",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"77",X"77",X"77",X"77",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"77",X"77",X"77",X"77",X"FF",X"FF",X"FF",X"FF",
		X"9F",X"66",X"FF",X"FF",X"FF",X"66",X"FF",X"FF",X"9F",X"66",X"FF",X"FF",X"9F",X"66",X"FF",X"FF",
		X"9F",X"66",X"FF",X"FF",X"CF",X"66",X"FF",X"FF",X"FF",X"6E",X"FF",X"FF",X"AF",X"6E",X"FF",X"FF",
		X"66",X"60",X"FF",X"FF",X"F6",X"EF",X"FF",X"FF",X"C7",X"EF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"66",X"FF",X"FF",X"FF",X"66",X"FF",X"FF",X"FF",X"66",X"FF",X"FF",X"FF",
		X"9F",X"99",X"66",X"FF",X"9F",X"99",X"66",X"FF",X"9F",X"99",X"66",X"FF",X"9F",X"9F",X"66",X"FF",
		X"9F",X"9F",X"6D",X"FF",X"9F",X"9F",X"6D",X"FF",X"9F",X"F6",X"6F",X"FF",X"9F",X"F6",X"DF",X"FF",
		X"9F",X"F6",X"DF",X"FF",X"9F",X"66",X"FF",X"FF",X"9F",X"66",X"FF",X"FF",X"9F",X"66",X"FF",X"FF",
		X"9F",X"66",X"FF",X"FF",X"9F",X"66",X"FF",X"FF",X"9F",X"66",X"FF",X"FF",X"9F",X"66",X"FF",X"FF",
		X"C4",X"44",X"44",X"7F",X"4C",X"44",X"44",X"7F",X"44",X"44",X"44",X"7F",X"C4",X"44",X"44",X"7F",
		X"4C",X"44",X"44",X"7F",X"CC",X"CC",X"CC",X"7F",X"99",X"99",X"99",X"7F",X"88",X"88",X"88",X"7F",
		X"88",X"88",X"88",X"7F",X"88",X"88",X"88",X"7F",X"88",X"88",X"88",X"7F",X"FF",X"FF",X"FF",X"7F",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"FF",X"FF",X"FF",X"FF",X"77",X"77",X"77",X"7F",X"CC",X"CC",X"CC",X"7F",X"CC",X"CC",X"CC",X"7F",
		X"CC",X"CC",X"CC",X"7F",X"CC",X"CC",X"CC",X"7F",X"44",X"44",X"44",X"7F",X"44",X"44",X"44",X"7F",
		X"C4",X"44",X"44",X"7F",X"4C",X"44",X"44",X"7F",X"C4",X"44",X"44",X"7F",X"4C",X"44",X"4C",X"7F",
		X"44",X"44",X"44",X"7F",X"44",X"44",X"C4",X"7F",X"44",X"44",X"4C",X"7F",X"44",X"44",X"44",X"7F",
		X"7F",X"22",X"22",X"F9",X"7F",X"22",X"22",X"FF",X"7F",X"22",X"22",X"77",X"7F",X"C2",X"22",X"77",
		X"9F",X"CC",X"C2",X"97",X"FF",X"EE",X"EE",X"F7",X"99",X"77",X"79",X"F7",X"77",X"77",X"77",X"F7",
		X"FF",X"22",X"22",X"F7",X"7F",X"22",X"22",X"77",X"7F",X"22",X"22",X"77",X"7F",X"22",X"22",X"77",
		X"7F",X"22",X"2E",X"99",X"7F",X"22",X"2E",X"FF",X"7F",X"22",X"22",X"F7",X"7F",X"22",X"22",X"F7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",
		X"FF",X"FF",X"DF",X"FF",X"FD",X"FF",X"DD",X"AA",X"DF",X"EF",X"FD",X"EE",X"FF",X"EF",X"FF",X"FF",
		X"FF",X"EF",X"FF",X"FF",X"FF",X"EF",X"FF",X"FF",X"FF",X"EF",X"FF",X"FF",X"FF",X"EF",X"FF",X"FF",
		X"AF",X"FF",X"FF",X"FF",X"AF",X"FA",X"FF",X"FF",X"FF",X"FA",X"FA",X"FF",X"FF",X"FA",X"FA",X"FF",
		X"AA",X"CA",X"CC",X"CC",X"77",X"7F",X"22",X"22",X"77",X"7F",X"22",X"22",X"77",X"7F",X"22",X"22",
		X"77",X"7F",X"22",X"2C",X"77",X"7F",X"22",X"2C",X"77",X"7F",X"CC",X"2C",X"AA",X"AA",X"C2",X"AA",
		X"88",X"9F",X"C2",X"66",X"77",X"8F",X"C2",X"88",X"77",X"8F",X"CC",X"88",X"77",X"8F",X"2C",X"88",
		X"77",X"8F",X"DE",X"88",X"77",X"8F",X"AE",X"88",X"FF",X"7F",X"CC",X"77",X"66",X"66",X"66",X"66",
		X"EF",X"EF",X"FA",X"EF",X"FA",X"AF",X"FA",X"EF",X"FE",X"EF",X"FA",X"EF",X"CE",X"EF",X"FA",X"FF",
		X"FC",X"F6",X"FA",X"FF",X"CF",X"C6",X"FA",X"F6",X"FC",X"F6",X"FF",X"F8",X"CF",X"F9",X"FF",X"FF",
		X"EA",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"E9",X"AE",X"AA",X"A2",X"C9",X"AA",X"AA",X"EC",X"CC",
		X"AA",X"AA",X"CC",X"CC",X"AA",X"2A",X"CC",X"CC",X"2E",X"E2",X"22",X"C6",X"66",X"66",X"66",X"66",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"FF",X"FF",X"FA",X"FF",X"FF",X"FF",X"EA",X"EF",X"FF",X"FF",X"EA",X"EF",X"EE",X"FF",
		X"EA",X"EF",X"AA",X"FF",X"FA",X"FA",X"EA",X"FF",X"EA",X"EF",X"EA",X"FF",X"EA",X"EF",X"AF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"FF",X"FF",X"FF",X"FE",
		X"88",X"AA",X"FF",X"FE",X"88",X"AA",X"FF",X"FE",X"88",X"7A",X"FF",X"EE",X"FF",X"FA",X"FF",X"FE",
		X"CC",X"CC",X"CC",X"AA",X"CC",X"CC",X"CC",X"AA",X"C2",X"CC",X"22",X"AA",X"22",X"CC",X"22",X"AE",
		X"22",X"CC",X"22",X"EE",X"C2",X"22",X"22",X"EE",X"C2",X"22",X"22",X"EE",X"CC",X"2C",X"CC",X"EE",
		X"CC",X"2C",X"CC",X"EE",X"C2",X"22",X"22",X"EE",X"99",X"99",X"99",X"EE",X"77",X"77",X"77",X"EE",
		X"99",X"99",X"99",X"EE",X"77",X"77",X"77",X"EA",X"77",X"77",X"77",X"AC",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"CC",X"C7",X"66",X"66",X"CC",X"C7",X"66",X"66",X"CC",X"76",
		X"66",X"67",X"EE",X"76",X"EE",X"EE",X"FF",X"EE",X"EE",X"EE",X"FF",X"EE",X"F9",X"FE",X"EE",X"99",
		X"99",X"FF",X"FF",X"99",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"96",X"FF",X"5D",X"DF",X"FF",
		X"FF",X"55",X"FF",X"FF",X"FF",X"DD",X"AF",X"FF",X"FF",X"5D",X"AF",X"FF",X"FF",X"AA",X"FF",X"FF",
		X"66",X"66",X"66",X"66",X"66",X"66",X"CC",X"C7",X"66",X"66",X"CC",X"C7",X"66",X"66",X"CC",X"76",
		X"66",X"67",X"EE",X"76",X"EE",X"5E",X"FF",X"EE",X"EE",X"E5",X"FF",X"EE",X"F5",X"EE",X"EE",X"99",
		X"C3",X"53",X"FF",X"99",X"33",X"5E",X"FF",X"FF",X"F5",X"EE",X"FF",X"96",X"FF",X"E5",X"FF",X"FF",
		X"FF",X"5E",X"EF",X"FF",X"FF",X"AA",X"EF",X"FF",X"FF",X"AA",X"FF",X"FF",X"FF",X"AA",X"FF",X"FF",
		X"66",X"D5",X"66",X"66",X"66",X"DD",X"5C",X"C7",X"66",X"D5",X"3C",X"C7",X"66",X"DD",X"3C",X"76",
		X"66",X"DD",X"EB",X"76",X"EB",X"FF",X"FF",X"EE",X"EE",X"EE",X"FB",X"EE",X"FF",X"99",X"BE",X"99",
		X"F8",X"77",X"FF",X"99",X"FF",X"17",X"FF",X"FF",X"FF",X"77",X"FF",X"96",X"FF",X"F6",X"FF",X"FF",
		X"FF",X"FF",X"AF",X"FF",X"FF",X"FF",X"AF",X"FF",X"FF",X"66",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"CC",X"CC",X"CC",X"CC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"CC",X"CC",X"CC",X"CC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"EE",X"FF",X"FF",X"EE",X"FF",X"FF",X"FF",X"FF",X"EF",X"FE",X"EE",X"EF",X"DE",X"ED",
		X"DD",X"E7",X"EE",X"DD",X"DD",X"7E",X"DD",X"DD",X"DD",X"67",X"DD",X"DD",X"DD",X"2E",X"DD",X"DD",
		X"DA",X"FD",X"FA",X"AF",X"DA",X"FF",X"FA",X"AF",X"DA",X"FF",X"FA",X"FF",X"DA",X"FF",X"AF",X"FF",
		X"AA",X"FF",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"DD",X"D7",X"7C",X"CC",X"DD",X"77",X"7C",X"CC",X"DD",X"C7",X"7C",X"CC",X"77",X"C7",X"7C",X"CC",
		X"CC",X"C7",X"7C",X"CC",X"77",X"C7",X"7C",X"CC",X"77",X"C7",X"7C",X"CC",X"77",X"C7",X"7C",X"CC",
		X"77",X"C7",X"7C",X"CC",X"77",X"77",X"7C",X"CC",X"CC",X"77",X"7C",X"CC",X"CC",X"77",X"7C",X"CC",
		X"CC",X"77",X"7C",X"CC",X"CC",X"77",X"7C",X"CC",X"CC",X"77",X"7C",X"CC",X"CC",X"77",X"7C",X"CC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FF",X"FF",X"EF",X"AE",
		X"FF",X"FF",X"EE",X"EE",X"FF",X"FE",X"DD",X"EA",X"FF",X"EE",X"DD",X"AF",X"EE",X"FF",X"DD",X"AF",
		X"DD",X"ED",X"AA",X"AF",X"DE",X"DD",X"AF",X"AF",X"EE",X"DD",X"FA",X"AF",X"DD",X"DD",X"FA",X"AF",
		X"DD",X"DD",X"FA",X"AF",X"DA",X"AD",X"FA",X"AF",X"DA",X"FD",X"FA",X"AF",X"DA",X"FD",X"FA",X"AF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"7C",
		X"FF",X"FF",X"FF",X"9C",X"FF",X"FF",X"FF",X"8C",X"FF",X"FF",X"FF",X"8C",X"FF",X"FF",X"FF",X"8C",
		X"FF",X"FF",X"F8",X"8C",X"FF",X"FF",X"87",X"8C",X"FF",X"FF",X"8C",X"8C",X"FF",X"FF",X"8C",X"8C",
		X"FF",X"FE",X"8C",X"8C",X"FF",X"ED",X"7C",X"8C",X"FE",X"DE",X"7C",X"8C",X"DD",X"D7",X"7C",X"8C",
		X"C7",X"77",X"7C",X"C7",X"C7",X"77",X"7C",X"C7",X"C7",X"77",X"7C",X"C7",X"C7",X"77",X"7C",X"C7",
		X"C7",X"77",X"7C",X"C7",X"C7",X"77",X"76",X"C7",X"C7",X"77",X"76",X"C7",X"C7",X"77",X"F9",X"C7",
		X"77",X"87",X"F9",X"C7",X"C7",X"C7",X"F9",X"C7",X"C7",X"C7",X"F9",X"77",X"C7",X"C7",X"F9",X"77",
		X"AA",X"C7",X"F9",X"77",X"AA",X"AA",X"F9",X"77",X"AA",X"AA",X"AA",X"77",X"AA",X"AA",X"AA",X"AA",
		X"11",X"11",X"11",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FB",X"BF",X"17",X"FB",X"FB",X"FB",X"17",
		X"FB",X"FB",X"BF",X"17",X"BB",X"FB",X"FB",X"17",X"FF",X"FF",X"FF",X"77",X"11",X"11",X"11",X"88",
		X"FF",X"FF",X"88",X"88",X"FF",X"FF",X"88",X"88",X"FF",X"FF",X"88",X"87",X"F1",X"FF",X"88",X"77",
		X"1F",X"F8",X"88",X"77",X"1F",X"88",X"88",X"77",X"11",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"FF",X"11",X"11",X"11",X"7F",X"FF",X"FF",X"FF",X"71",X"BB",X"FF",X"FB",X"71",X"FF",X"BF",X"FB",
		X"71",X"FF",X"BF",X"FB",X"71",X"BB",X"FF",X"FB",X"77",X"FF",X"FF",X"FF",X"77",X"11",X"11",X"FF",
		X"77",X"FF",X"F1",X"1F",X"77",X"88",X"81",X"1F",X"77",X"88",X"81",X"FF",X"77",X"88",X"71",X"1F",
		X"78",X"88",X"71",X"1F",X"88",X"88",X"71",X"1F",X"99",X"99",X"71",X"FF",X"99",X"99",X"78",X"88",
		X"7F",X"22",X"22",X"66",X"7F",X"22",X"22",X"FF",X"7F",X"22",X"22",X"77",X"7F",X"22",X"22",X"77",
		X"7F",X"22",X"22",X"77",X"7F",X"22",X"22",X"77",X"7F",X"22",X"22",X"77",X"7F",X"CC",X"CC",X"66",
		X"77",X"88",X"88",X"66",X"7F",X"22",X"22",X"FF",X"7F",X"22",X"22",X"77",X"7F",X"22",X"22",X"77",
		X"7F",X"22",X"22",X"77",X"7F",X"22",X"22",X"77",X"7F",X"22",X"22",X"77",X"7F",X"22",X"22",X"66",
		X"FF",X"96",X"88",X"98",X"FF",X"96",X"88",X"98",X"FF",X"96",X"88",X"98",X"A2",X"AA",X"A2",X"AA",
		X"E2",X"2E",X"22",X"2E",X"EE",X"EE",X"EE",X"EE",X"11",X"E1",X"1E",X"EE",X"1E",X"E1",X"EE",X"EE",
		X"11",X"E1",X"EE",X"EE",X"1E",X"E1",X"EE",X"EE",X"EE",X"E1",X"EE",X"EE",X"33",X"11",X"1E",X"EE",
		X"3E",X"EE",X"EE",X"EE",X"33",X"AA",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"77",X"77",X"77",X"77",
		X"FF",X"99",X"FF",X"FF",X"79",X"55",X"99",X"FF",X"75",X"55",X"59",X"FF",X"75",X"55",X"59",X"FF",
		X"75",X"55",X"59",X"FF",X"75",X"55",X"59",X"FF",X"79",X"88",X"59",X"FF",X"79",X"88",X"69",X"FF",
		X"79",X"55",X"69",X"FF",X"75",X"55",X"59",X"FF",X"75",X"55",X"59",X"FF",X"75",X"55",X"59",X"FF",
		X"75",X"55",X"59",X"FF",X"75",X"55",X"59",X"FF",X"89",X"88",X"59",X"FF",X"89",X"88",X"69",X"FF",
		X"8A",X"8A",X"8A",X"FA",X"8A",X"8A",X"8A",X"FF",X"8A",X"8A",X"8A",X"FF",X"8A",X"8A",X"8A",X"FE",
		X"8A",X"8A",X"8A",X"EE",X"8A",X"8A",X"8A",X"EE",X"8A",X"8A",X"8A",X"EE",X"8A",X"8A",X"8A",X"EF",
		X"8A",X"8A",X"8A",X"FE",X"8A",X"8A",X"8A",X"EE",X"8A",X"8A",X"8A",X"EE",X"8A",X"8A",X"8A",X"EE",
		X"8A",X"8A",X"8A",X"EA",X"8A",X"8A",X"8A",X"AA",X"77",X"77",X"77",X"AC",X"66",X"66",X"66",X"66",
		X"76",X"EA",X"8A",X"8A",X"AF",X"EA",X"8A",X"8A",X"AF",X"EA",X"8A",X"8A",X"AF",X"EA",X"8A",X"8A",
		X"AF",X"FA",X"9A",X"8A",X"AF",X"FF",X"9A",X"8A",X"AF",X"FF",X"9A",X"8A",X"AF",X"FF",X"9A",X"8A",
		X"AF",X"FF",X"9A",X"8A",X"AF",X"FF",X"9A",X"8A",X"AF",X"FF",X"8A",X"8A",X"AF",X"FF",X"8A",X"8A",
		X"A6",X"FF",X"8A",X"8A",X"66",X"FF",X"8A",X"8A",X"FF",X"F6",X"76",X"76",X"FF",X"66",X"66",X"66",
		X"77",X"FF",X"77",X"77",X"77",X"FF",X"99",X"99",X"77",X"FF",X"88",X"88",X"77",X"FF",X"7A",X"7A",
		X"77",X"FF",X"FA",X"7A",X"77",X"FF",X"7A",X"7A",X"77",X"FF",X"7A",X"7A",X"77",X"FF",X"88",X"88",
		X"77",X"FF",X"99",X"99",X"77",X"EF",X"88",X"88",X"77",X"ED",X"7A",X"7A",X"77",X"DD",X"7A",X"7A",
		X"77",X"DD",X"7A",X"8A",X"77",X"DA",X"8A",X"8A",X"77",X"DA",X"8A",X"8A",X"77",X"FA",X"8A",X"8A",
		X"77",X"77",X"77",X"77",X"99",X"99",X"99",X"99",X"77",X"88",X"88",X"77",X"99",X"99",X"99",X"99",
		X"77",X"88",X"88",X"77",X"99",X"99",X"99",X"99",X"77",X"88",X"88",X"88",X"99",X"99",X"FF",X"FF",
		X"99",X"99",X"F7",X"77",X"77",X"88",X"F7",X"77",X"FF",X"FF",X"F7",X"77",X"77",X"77",X"77",X"77",
		X"88",X"88",X"88",X"88",X"99",X"99",X"99",X"99",X"88",X"88",X"88",X"88",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"87",X"8F",X"FF",X"7F",X"87",X"8F",X"FF",X"7F",X"87",X"8F",X"FF",X"7F",X"8A",X"7F",X"FF",
		X"7F",X"8A",X"7F",X"FF",X"7F",X"AA",X"7F",X"FF",X"7F",X"AA",X"7F",X"FF",X"7F",X"A8",X"8F",X"FF",
		X"7F",X"A8",X"8F",X"FF",X"7F",X"88",X"8F",X"FF",X"7F",X"88",X"8F",X"FF",X"7F",X"88",X"8F",X"FF",
		X"7F",X"88",X"8F",X"FF",X"7F",X"88",X"8F",X"FF",X"7F",X"88",X"8F",X"FF",X"7A",X"88",X"8F",X"FF",
		X"88",X"AA",X"AA",X"99",X"99",X"AC",X"AC",X"9D",X"99",X"AC",X"AC",X"9D",X"C6",X"AC",X"A2",X"97",
		X"CC",X"A2",X"A2",X"97",X"C6",X"E2",X"A2",X"97",X"66",X"E2",X"A2",X"97",X"C6",X"D2",X"A2",X"97",
		X"CC",X"D2",X"A2",X"97",X"99",X"D2",X"A2",X"96",X"99",X"D2",X"A2",X"97",X"77",X"DD",X"AA",X"99",
		X"99",X"CC",X"CC",X"99",X"99",X"CC",X"CC",X"99",X"88",X"CC",X"CC",X"77",X"66",X"66",X"66",X"66",
		X"8A",X"88",X"CA",X"FF",X"AA",X"88",X"2A",X"FF",X"AA",X"88",X"2A",X"FF",X"EF",X"88",X"2A",X"FF",
		X"EF",X"88",X"2A",X"FF",X"7F",X"88",X"2A",X"FF",X"7F",X"88",X"CA",X"FF",X"7F",X"88",X"CA",X"FF",
		X"7F",X"88",X"2A",X"FF",X"7F",X"88",X"AA",X"FF",X"7F",X"89",X"99",X"FF",X"7F",X"89",X"77",X"FF",
		X"7F",X"DD",X"7F",X"FF",X"7F",X"DD",X"EA",X"FF",X"7F",X"DD",X"DA",X"FF",X"7F",X"DD",X"DA",X"FF",
		X"FF",X"72",X"FE",X"2E",X"EE",X"72",X"EE",X"2E",X"77",X"77",X"7F",X"7F",X"77",X"72",X"8F",X"2F",
		X"77",X"72",X"8F",X"2F",X"77",X"77",X"8F",X"7F",X"78",X"72",X"8F",X"2F",X"88",X"72",X"9F",X"2F",
		X"88",X"77",X"9F",X"7F",X"89",X"72",X"9F",X"2F",X"99",X"72",X"9F",X"CF",X"99",X"77",X"9F",X"7F",
		X"99",X"7C",X"9F",X"CF",X"99",X"7C",X"9F",X"CF",X"99",X"77",X"9F",X"7F",X"99",X"7C",X"9F",X"CF",
		X"77",X"88",X"88",X"9F",X"AA",X"AC",X"FF",X"A8",X"CC",X"AC",X"FF",X"AA",X"CC",X"AC",X"77",X"AA",
		X"C2",X"A2",X"77",X"AA",X"C2",X"A2",X"77",X"AA",X"C2",X"A2",X"77",X"AA",X"C2",X"A2",X"77",X"AE",
		X"C2",X"A2",X"77",X"AE",X"C2",X"A2",X"77",X"AE",X"C2",X"A2",X"77",X"AE",X"C2",X"AC",X"77",X"AA",
		X"CC",X"A2",X"CC",X"AA",X"CC",X"AF",X"CC",X"AA",X"AA",X"CC",X"CC",X"AC",X"66",X"66",X"66",X"66",
		X"44",X"77",X"77",X"77",X"44",X"77",X"77",X"77",X"4F",X"70",X"77",X"77",X"44",X"77",X"77",X"77",
		X"44",X"77",X"77",X"77",X"4F",X"70",X"77",X"77",X"4F",X"70",X"77",X"77",X"7F",X"77",X"77",X"77",
		X"4F",X"77",X"77",X"77",X"44",X"70",X"77",X"77",X"44",X"77",X"77",X"77",X"4F",X"77",X"77",X"77",
		X"4F",X"70",X"77",X"77",X"4F",X"70",X"77",X"77",X"FF",X"F0",X"FF",X"FF",X"7F",X"77",X"77",X"77",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"44",X"FF",X"FF",X"F4",X"4F",X"4F",
		X"FF",X"F4",X"44",X"4F",X"FF",X"F4",X"4F",X"4F",X"FF",X"F4",X"44",X"4F",X"FF",X"F4",X"FF",X"FF",
		X"FF",X"44",X"F1",X"11",X"FF",X"FF",X"FF",X"1F",X"FF",X"FF",X"FF",X"11",X"FF",X"FF",X"FF",X"1F",
		X"88",X"88",X"81",X"11",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",
		X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"C7",X"FF",X"FF",X"FF",X"C7",X"FF",X"FF",X"FF",
		X"C7",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",
		X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DD",X"DD",X"DD",
		X"DD",X"55",X"55",X"D5",X"99",X"CC",X"CC",X"AC",X"99",X"CC",X"CC",X"AC",X"99",X"C5",X"5C",X"A5",
		X"99",X"C5",X"5C",X"A5",X"99",X"C5",X"5C",X"A5",X"99",X"C5",X"5C",X"A5",X"99",X"CC",X"5C",X"A5",
		X"99",X"CC",X"5C",X"A5",X"99",X"CC",X"5C",X"A5",X"88",X"88",X"88",X"88",X"77",X"EE",X"EE",X"EE",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"77",X"77",X"77",X"77",X"45",X"45",X"45",X"47",X"45",X"45",X"45",X"47",X"45",X"45",X"45",X"11",
		X"53",X"53",X"53",X"57",X"53",X"53",X"53",X"00",X"53",X"53",X"53",X"57",X"34",X"34",X"34",X"BB",
		X"34",X"34",X"34",X"37",X"34",X"34",X"34",X"37",X"77",X"77",X"77",X"77",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"7F",X"F7",X"F7",X"7F",X"7F",X"F7",X"F7",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"77",X"77",X"77",X"77",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",
		X"53",X"53",X"53",X"53",X"53",X"53",X"53",X"53",X"53",X"53",X"53",X"53",X"34",X"34",X"34",X"34",
		X"34",X"34",X"34",X"34",X"34",X"34",X"34",X"34",X"77",X"77",X"77",X"77",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"22",X"22",X"66",X"7F",X"22",X"22",X"FF",X"7F",X"0C",X"04",X"77",X"7F",X"C0",X"CC",X"77",
		X"7F",X"2C",X"22",X"77",X"CC",X"CC",X"22",X"77",X"00",X"00",X"22",X"77",X"7F",X"CC",X"CC",X"66",
		X"77",X"88",X"88",X"66",X"7F",X"24",X"2C",X"FF",X"4F",X"4C",X"C4",X"77",X"4F",X"4C",X"C4",X"77",
		X"7F",X"4C",X"2C",X"77",X"4F",X"4C",X"CC",X"77",X"7F",X"C2",X"44",X"77",X"7F",X"22",X"CC",X"66",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"4F",X"4F",X"FF",X"FF",X"4F",X"FF",X"4F",X"FF",
		X"44",X"FF",X"FF",X"FF",X"4F",X"FF",X"FF",X"FF",X"4F",X"4F",X"44",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"F4",X"FF",X"FF",X"1F",X"FF",X"FF",X"FF",X"1F",X"FF",X"FF",X"FF",X"1F",X"FF",X"FF",X"FF",
		X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"99",X"99",X"98",X"FF",X"98",X"98",X"89",X"FF",X"89",X"89",X"99",X"FF",
		X"99",X"99",X"97",X"FF",X"99",X"9F",X"87",X"FF",X"F9",X"F8",X"CA",X"FF",X"8F",X"F8",X"2A",X"FF",
		X"99",X"C8",X"2A",X"FF",X"99",X"F8",X"2A",X"FF",X"99",X"C7",X"2A",X"FF",X"99",X"77",X"CA",X"FF",
		X"99",X"77",X"2A",X"FF",X"99",X"78",X"2A",X"FF",X"99",X"77",X"FA",X"FF",X"9F",X"77",X"99",X"FF",
		X"88",X"CC",X"CC",X"AA",X"88",X"CC",X"CC",X"AA",X"88",X"22",X"22",X"AA",X"99",X"2C",X"CC",X"AE",
		X"99",X"CC",X"CC",X"EE",X"99",X"2C",X"CC",X"EE",X"99",X"CC",X"2C",X"EE",X"99",X"CC",X"2C",X"EE",
		X"99",X"C2",X"CC",X"EE",X"99",X"CC",X"CC",X"EE",X"99",X"C2",X"CC",X"EE",X"99",X"CC",X"CC",X"EE",
		X"99",X"CC",X"CC",X"EE",X"99",X"99",X"99",X"EA",X"99",X"77",X"77",X"AC",X"66",X"66",X"66",X"66",
		X"55",X"55",X"77",X"F7",X"55",X"55",X"77",X"F7",X"7F",X"F7",X"77",X"FF",X"7F",X"55",X"55",X"F5",
		X"7F",X"55",X"5F",X"5F",X"7F",X"55",X"5F",X"F5",X"7F",X"F5",X"5F",X"F7",X"7F",X"FF",X"FF",X"FF",
		X"7F",X"77",X"BB",X"BB",X"7F",X"77",X"BB",X"BB",X"7F",X"77",X"F3",X"FF",X"7F",X"77",X"33",X"33",
		X"7F",X"77",X"33",X"33",X"7F",X"77",X"F4",X"FA",X"7F",X"77",X"44",X"FF",X"7F",X"77",X"44",X"FA",
		X"77",X"F5",X"77",X"F7",X"5F",X"F5",X"77",X"F7",X"FF",X"F5",X"77",X"F7",X"5F",X"F5",X"77",X"55",
		X"5F",X"F5",X"F7",X"FF",X"5F",X"F5",X"F7",X"5F",X"5F",X"55",X"5F",X"FF",X"FC",X"FF",X"AA",X"FF",
		X"BB",X"BB",X"FF",X"FF",X"BB",X"BB",X"FF",X"5F",X"F3",X"33",X"F7",X"5F",X"73",X"33",X"F7",X"55",
		X"73",X"33",X"F7",X"F7",X"74",X"44",X"F7",X"F7",X"74",X"44",X"F7",X"F7",X"74",X"44",X"F7",X"F7",
		X"FF",X"FF",X"FF",X"FC",X"99",X"99",X"FF",X"9C",X"77",X"FF",X"FF",X"FC",X"88",X"99",X"99",X"88",
		X"88",X"99",X"99",X"98",X"8E",X"99",X"88",X"78",X"9E",X"89",X"98",X"88",X"99",X"8F",X"99",X"88",
		X"99",X"98",X"99",X"88",X"99",X"98",X"77",X"99",X"99",X"FF",X"99",X"9C",X"FF",X"8F",X"99",X"FC",
		X"99",X"88",X"99",X"88",X"99",X"88",X"99",X"88",X"77",X"C8",X"77",X"78",X"77",X"99",X"77",X"79",
		X"FF",X"66",X"66",X"66",X"FF",X"66",X"66",X"66",X"FF",X"66",X"66",X"66",X"FF",X"88",X"88",X"88",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"8F",X"66",X"66",X"66",X"FF",X"88",X"88",X"88",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"89",X"88",X"69",X"FF",X"89",X"88",X"69",X"FF",X"89",X"88",X"69",X"FF",X"A2",X"AA",X"A2",X"AA",
		X"22",X"2E",X"22",X"E2",X"EE",X"EE",X"EE",X"EE",X"EE",X"E1",X"E1",X"EE",X"EE",X"EE",X"E1",X"E1",
		X"EE",X"EE",X"E1",X"E1",X"EE",X"EE",X"E1",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"E1",X"3E",X"3E",
		X"EE",X"EE",X"33",X"3E",X"AA",X"AA",X"3A",X"3A",X"FF",X"FF",X"FF",X"FF",X"77",X"77",X"77",X"77",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"88",X"88",X"88",X"88",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"89",X"88",X"69",X"FF",X"89",X"88",X"69",X"FF",X"89",X"88",X"69",X"FF",X"89",X"88",X"69",X"FF",
		X"89",X"88",X"69",X"FF",X"89",X"88",X"69",X"FF",X"89",X"88",X"69",X"FF",X"89",X"88",X"69",X"FF",
		X"89",X"88",X"69",X"FF",X"ED",X"88",X"69",X"FF",X"89",X"AE",X"DA",X"FF",X"89",X"77",X"78",X"FF",
		X"89",X"77",X"88",X"FF",X"89",X"77",X"88",X"FC",X"89",X"CC",X"CC",X"CC",X"66",X"66",X"66",X"66",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",
		X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"C7",X"FF",X"FF",X"FF",X"C7",X"FF",X"FF",X"FF",
		X"C7",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",
		X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"2F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"99",X"FF",X"FF",X"FF",X"55",X"FF",X"FF",X"FF",X"55",
		X"FF",X"FF",X"FF",X"55",X"FF",X"FF",X"FF",X"99",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"99",
		X"7A",X"77",X"DD",X"FF",X"A7",X"7A",X"FF",X"FF",X"FF",X"7A",X"FF",X"AF",X"FC",X"7A",X"FF",X"FF",
		X"FC",X"CC",X"FF",X"FF",X"99",X"99",X"FF",X"6F",X"88",X"88",X"FF",X"CF",X"99",X"99",X"9F",X"CF",
		X"88",X"88",X"9F",X"99",X"88",X"88",X"9F",X"88",X"77",X"88",X"9F",X"88",X"77",X"88",X"9F",X"88",
		X"77",X"88",X"9F",X"88",X"77",X"88",X"9F",X"88",X"77",X"88",X"9F",X"77",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"9F",X"FF",X"FF",X"FF",X"79",X"F0",X"00",X"09",X"97",X"F0",X"0F",X"90",
		X"09",X"F0",X"00",X"70",X"07",X"F0",X"0F",X"90",X"70",X"F0",X"00",X"09",X"97",X"9F",X"FF",X"97",
		X"99",X"33",X"39",X"79",X"F9",X"37",X"37",X"99",X"FF",X"33",X"39",X"9F",X"FF",X"99",X"99",X"F7",
		X"FF",X"FF",X"FF",X"F8",X"99",X"99",X"99",X"99",X"88",X"88",X"88",X"88",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"88",X"88",X"88",X"88",X"8A",X"CC",X"8F",X"88",X"AA",X"CC",X"F8",X"77",X"FF",X"FF",X"F7",
		X"77",X"EA",X"CC",X"F7",X"77",X"EE",X"CC",X"F7",X"77",X"EE",X"CC",X"F7",X"77",X"EE",X"22",X"F7",
		X"77",X"EE",X"22",X"F7",X"77",X"EE",X"22",X"F7",X"77",X"EE",X"22",X"F7",X"77",X"EE",X"22",X"F7",
		X"77",X"EE",X"22",X"F7",X"77",X"EE",X"22",X"F7",X"77",X"EE",X"22",X"F7",X"77",X"AE",X"22",X"F7",
		X"88",X"88",X"88",X"88",X"88",X"88",X"A2",X"CC",X"8F",X"8F",X"22",X"CC",X"F7",X"F7",X"FF",X"FF",
		X"F7",X"F7",X"CC",X"CE",X"F7",X"F7",X"CC",X"2E",X"F7",X"F7",X"CC",X"2A",X"F7",X"F7",X"CC",X"2A",
		X"F7",X"F7",X"CC",X"2A",X"F7",X"F7",X"CC",X"2A",X"F7",X"F7",X"C2",X"2A",X"F7",X"F7",X"C2",X"2A",
		X"F7",X"F7",X"22",X"2A",X"F7",X"F7",X"22",X"2F",X"F7",X"F7",X"22",X"2F",X"F7",X"F7",X"22",X"2F",
		X"78",X"77",X"67",X"FA",X"77",X"77",X"67",X"FA",X"87",X"87",X"67",X"FA",X"88",X"87",X"67",X"FA",
		X"88",X"87",X"67",X"FA",X"88",X"87",X"67",X"FA",X"88",X"88",X"67",X"FA",X"88",X"87",X"67",X"FA",
		X"88",X"87",X"67",X"FA",X"88",X"87",X"67",X"FA",X"88",X"87",X"67",X"FA",X"88",X"77",X"67",X"FA",
		X"FF",X"77",X"67",X"FA",X"AA",X"77",X"67",X"FA",X"AA",X"FF",X"67",X"F6",X"AA",X"AA",X"67",X"66",
		X"AA",X"AA",X"6A",X"AA",X"77",X"77",X"66",X"77",X"A7",X"A7",X"66",X"EE",X"FA",X"FA",X"66",X"FF",
		X"FA",X"CA",X"66",X"CC",X"FA",X"CA",X"66",X"CC",X"FA",X"CA",X"F6",X"CC",X"FA",X"CA",X"66",X"CC",
		X"CC",X"2A",X"66",X"22",X"2C",X"2A",X"66",X"22",X"2C",X"2A",X"66",X"22",X"AC",X"2A",X"66",X"FF",
		X"FC",X"DE",X"86",X"FF",X"CC",X"88",X"68",X"EE",X"FF",X"77",X"67",X"77",X"78",X"77",X"67",X"9F",
		X"FF",X"FF",X"6F",X"FF",X"FF",X"FF",X"69",X"6F",X"FF",X"FA",X"C9",X"77",X"FF",X"A8",X"CE",X"77",
		X"FA",X"88",X"97",X"77",X"A8",X"88",X"77",X"FF",X"88",X"AA",X"77",X"88",X"8F",X"FC",X"7F",X"88",
		X"AF",X"FC",X"F8",X"88",X"A2",X"FC",X"88",X"88",X"A2",X"F2",X"88",X"88",X"A2",X"F2",X"78",X"88",
		X"68",X"F2",X"77",X"88",X"68",X"FF",X"77",X"88",X"68",X"FF",X"17",X"88",X"77",X"77",X"77",X"77",
		X"CF",X"FF",X"FF",X"77",X"11",X"F1",X"11",X"F1",X"F1",X"81",X"DD",X"1F",X"F1",X"F1",X"1D",X"F1",
		X"F1",X"F1",X"AA",X"F7",X"F1",X"11",X"11",X"11",X"88",X"88",X"88",X"7F",X"AA",X"71",X"18",X"7F",
		X"9A",X"71",X"18",X"7F",X"98",X"F1",X"18",X"7F",X"98",X"F1",X"18",X"7F",X"9A",X"F1",X"11",X"7A",
		X"97",X"88",X"FF",X"7A",X"CC",X"CC",X"AA",X"7A",X"CC",X"CC",X"97",X"CC",X"CC",X"CC",X"99",X"CC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"FF",
		X"FF",X"FF",X"FC",X"CC",X"FF",X"FF",X"FC",X"CF",X"FF",X"FF",X"FC",X"CF",X"FF",X"FF",X"77",X"77",
		X"79",X"FF",X"FF",X"FC",X"79",X"DF",X"AA",X"FF",X"79",X"DD",X"AF",X"AF",X"79",X"DA",X"AF",X"FF",
		X"79",X"FF",X"AF",X"6F",X"79",X"FF",X"FF",X"99",X"79",X"FF",X"FF",X"77",X"79",X"FF",X"FF",X"77",
		X"79",X"FF",X"FF",X"77",X"79",X"FF",X"66",X"77",X"78",X"A6",X"67",X"77",X"78",X"67",X"77",X"77",
		X"78",X"7F",X"77",X"7F",X"77",X"22",X"77",X"FF",X"77",X"FC",X"FF",X"FC",X"77",X"CC",X"CC",X"CC",
		X"FF",X"FF",X"AA",X"AA",X"FF",X"FF",X"FC",X"CC",X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"CC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"FF",X"FF",X"FF",X"CF",X"FF",X"FF",X"CC",X"CC",
		X"F7",X"FF",X"CF",X"CC",X"F7",X"FF",X"CF",X"CF",X"F7",X"FF",X"CF",X"CF",X"F8",X"FF",X"CF",X"CF",
		X"F6",X"9F",X"CC",X"CC",X"F9",X"FF",X"FF",X"FF",X"79",X"FF",X"FF",X"CC",X"79",X"FF",X"FF",X"CF",
		X"AA",X"AA",X"6A",X"CC",X"AA",X"AA",X"AA",X"CC",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"AA",
		X"AA",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AD",X"EA",X"AA",X"AA",X"AF",X"AA",X"AA",X"AA",
		X"AA",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"AA",X"AA",X"AA",X"CE",X"AA",X"AE",
		X"AA",X"EA",X"DA",X"AA",X"AA",X"AA",X"ED",X"AA",X"CC",X"FC",X"EE",X"66",X"CC",X"CC",X"CF",X"C6",
		X"77",X"CC",X"CC",X"CC",X"77",X"CC",X"CC",X"CC",X"77",X"C6",X"66",X"AA",X"77",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"22",X"CC",X"AA",X"CC",X"CC",X"CC",X"AA",X"C8",X"CC",X"CA",X"AA",X"EE",X"CC",X"AA",
		X"AA",X"EE",X"CA",X"AA",X"AA",X"AA",X"AA",X"AA",X"CA",X"AA",X"AA",X"EE",X"CA",X"AA",X"AA",X"EF",
		X"FC",X"AA",X"AA",X"EE",X"FC",X"AA",X"AA",X"AA",X"FF",X"CE",X"66",X"6C",X"FF",X"CC",X"6F",X"6C",
		X"CC",X"CC",X"99",X"CC",X"CC",X"CC",X"99",X"CC",X"FF",X"FF",X"99",X"CC",X"FF",X"CC",X"77",X"AA",
		X"AC",X"CC",X"CC",X"AA",X"AA",X"CC",X"CC",X"AA",X"CA",X"AC",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EC",X"AA",X"AA",X"AA",X"AC",
		X"DD",X"AA",X"AA",X"6F",X"DA",X"AA",X"DD",X"6F",X"CC",X"CC",X"EC",X"FF",X"CC",X"CC",X"CC",X"FF",
		X"F7",X"77",X"FF",X"F1",X"F7",X"70",X"71",X"1F",X"F7",X"70",X"71",X"1F",X"87",X"70",X"71",X"1F",
		X"87",X"70",X"71",X"1F",X"87",X"70",X"7F",X"F1",X"87",X"70",X"7F",X"FF",X"87",X"70",X"74",X"4F",
		X"87",X"70",X"4F",X"FF",X"87",X"70",X"74",X"FF",X"87",X"70",X"7F",X"FF",X"87",X"70",X"44",X"88",
		X"87",X"70",X"77",X"70",X"87",X"70",X"77",X"70",X"87",X"70",X"77",X"70",X"69",X"2F",X"22",X"9F",
		X"FF",X"FF",X"F9",X"FF",X"FF",X"FF",X"97",X"6F",X"FF",X"FA",X"67",X"77",X"FF",X"A8",X"67",X"77",
		X"FA",X"88",X"97",X"77",X"A8",X"88",X"7C",X"FF",X"88",X"AA",X"77",X"88",X"8F",X"FC",X"7F",X"88",
		X"AF",X"FC",X"F8",X"88",X"A2",X"FC",X"88",X"88",X"A2",X"F2",X"88",X"88",X"A2",X"F2",X"78",X"88",
		X"68",X"F2",X"77",X"88",X"68",X"FF",X"77",X"88",X"68",X"FF",X"17",X"88",X"77",X"77",X"77",X"77",
		X"CF",X"FF",X"AA",X"AA",X"CF",X"FF",X"AA",X"AA",X"FF",X"FF",X"CA",X"AA",X"FF",X"FF",X"FC",X"CC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AD",X"DD",X"DA",X"AA",X"AD",X"DA",X"AF",X"AF",X"AD",X"EA",X"AF",X"AF",X"AD",X"DA",X"AF",X"AF",
		X"AD",X"AA",X"AF",X"FF",X"AA",X"FF",X"FA",X"FF",X"FF",X"FF",X"FA",X"AA",X"FF",X"FF",X"FF",X"FA",
		X"FF",X"FF",X"FF",X"FA",X"F2",X"FF",X"FF",X"FA",X"F7",X"FF",X"FF",X"FF",X"FC",X"AA",X"AA",X"AA",
		X"FF",X"AA",X"AA",X"AA",X"FF",X"FC",X"AA",X"AA",X"CF",X"FF",X"AA",X"AA",X"AC",X"FF",X"AA",X"AA",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"88",X"88",X"8F",X"88",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"99",X"99",X"FF",X"FF",X"77",X"77",X"FF",X"FF",
		X"88",X"88",X"FF",X"FF",X"88",X"89",X"FF",X"FF",X"88",X"98",X"FF",X"FF",X"88",X"88",X"FF",X"FF",
		X"87",X"88",X"FF",X"FF",X"7F",X"88",X"FF",X"FF",X"77",X"88",X"FF",X"FF",X"89",X"88",X"FF",X"FF",
		X"7F",X"DD",X"DA",X"FF",X"7F",X"DD",X"DA",X"FF",X"7F",X"DD",X"DA",X"FF",X"7F",X"DD",X"DA",X"FF",
		X"7F",X"DD",X"DA",X"FF",X"7F",X"ED",X"DA",X"DF",X"7F",X"ED",X"DA",X"DF",X"7F",X"ED",X"DA",X"FF",
		X"7A",X"ED",X"DA",X"FF",X"7F",X"ED",X"DA",X"FF",X"7F",X"EE",X"DA",X"FF",X"7F",X"EE",X"DA",X"FF",
		X"7F",X"EE",X"DA",X"FF",X"7F",X"EE",X"F6",X"FF",X"7F",X"EE",X"66",X"FF",X"7F",X"99",X"66",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",
		X"F7",X"EA",X"FF",X"FF",X"7F",X"DC",X"EA",X"FF",X"7F",X"DE",X"DA",X"FF",X"9F",X"DD",X"DA",X"FF",
		X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"F7",X"FF",X"FF",X"77",X"F7",X"FF",X"7F",X"77",X"F7",X"FF",
		X"77",X"EE",X"DE",X"99",X"9F",X"77",X"F7",X"97",X"9F",X"77",X"A7",X"99",X"9F",X"77",X"F7",X"99",
		X"9F",X"FF",X"F7",X"89",X"9F",X"FF",X"77",X"89",X"9F",X"FF",X"77",X"88",X"8F",X"FF",X"FF",X"8F",
		X"FF",X"FF",X"FF",X"87",X"FF",X"ED",X"AA",X"F8",X"7F",X"DD",X"AA",X"7F",X"8F",X"99",X"F9",X"F8",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"88",X"88",X"88",X"88",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"99",X"99",X"99",X"FF",X"77",X"77",X"7C",
		X"FF",X"88",X"88",X"8C",X"99",X"CC",X"8A",X"88",X"77",X"C8",X"88",X"88",X"88",X"A8",X"8F",X"88",
		X"88",X"88",X"FF",X"88",X"88",X"88",X"88",X"88",X"89",X"98",X"88",X"98",X"97",X"79",X"99",X"79",
		X"66",X"66",X"66",X"66",X"66",X"66",X"CC",X"C7",X"66",X"66",X"CC",X"C7",X"66",X"66",X"CC",X"76",
		X"66",X"67",X"EE",X"76",X"EE",X"EE",X"F1",X"EE",X"EE",X"EE",X"F8",X"EE",X"F9",X"FE",X"EE",X"99",
		X"99",X"FF",X"FF",X"99",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"96",X"FF",X"D5",X"FF",X"FF",
		X"FF",X"DD",X"5F",X"FF",X"FF",X"D5",X"DF",X"FF",X"FF",X"DD",X"FF",X"FF",X"FF",X"DD",X"FF",X"FF",
		X"66",X"FF",X"FF",X"FF",X"66",X"CF",X"FF",X"FF",X"66",X"FF",X"FF",X"FF",X"66",X"FF",X"FF",X"FF",
		X"6E",X"FF",X"FF",X"FF",X"EE",X"FF",X"FF",X"FF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"88",X"88",X"88",X"88",
		X"FF",X"FF",X"FF",X"FF",X"AC",X"FF",X"FF",X"FF",X"AC",X"99",X"99",X"99",X"AC",X"77",X"77",X"77",
		X"AC",X"88",X"88",X"88",X"AC",X"8A",X"88",X"88",X"AA",X"AA",X"88",X"FF",X"88",X"CC",X"88",X"88",
		X"8F",X"CC",X"88",X"88",X"88",X"88",X"88",X"88",X"99",X"88",X"99",X"89",X"77",X"99",X"77",X"97",
		X"9F",X"88",X"FF",X"FF",X"7F",X"88",X"FF",X"FF",X"7F",X"88",X"CF",X"FF",X"7F",X"88",X"CF",X"FF",
		X"7F",X"88",X"9F",X"FF",X"7F",X"88",X"9F",X"FF",X"7F",X"88",X"9F",X"FF",X"7F",X"88",X"9F",X"FF",
		X"7F",X"88",X"9F",X"FF",X"7F",X"88",X"9F",X"FF",X"7F",X"88",X"9F",X"FF",X"7F",X"88",X"DD",X"FF",
		X"7F",X"88",X"A8",X"FF",X"7F",X"88",X"AF",X"FF",X"7F",X"88",X"8F",X"FF",X"7F",X"88",X"8F",X"FF",
		X"F5",X"55",X"99",X"99",X"55",X"55",X"77",X"FF",X"55",X"FF",X"77",X"FF",X"55",X"77",X"77",X"FF",
		X"55",X"55",X"77",X"FF",X"55",X"FF",X"FF",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"5F",X"FF",X"FF",X"55",X"F5",X"F5",X"F5",X"FF",X"5F",X"5F",X"F5",
		X"FF",X"F2",X"F5",X"F5",X"55",X"57",X"F5",X"F5",X"FF",X"F5",X"55",X"F5",X"7F",X"5F",X"F5",X"FF",
		X"8A",X"85",X"8F",X"F5",X"AA",X"85",X"8F",X"F5",X"AA",X"85",X"85",X"F5",X"EF",X"85",X"8F",X"F5",
		X"EF",X"85",X"8F",X"F5",X"8F",X"88",X"8F",X"FF",X"8F",X"85",X"55",X"F5",X"8F",X"95",X"85",X"F5",
		X"8F",X"95",X"55",X"F5",X"8F",X"99",X"8F",X"FF",X"8F",X"99",X"8F",X"FF",X"8F",X"99",X"8F",X"FF",
		X"8F",X"DD",X"7F",X"FF",X"8F",X"DD",X"EA",X"FF",X"7F",X"DD",X"DA",X"FF",X"7F",X"DD",X"DA",X"FF",
		X"7F",X"DD",X"DA",X"FF",X"7E",X"DD",X"DA",X"FF",X"7F",X"DD",X"DA",X"FF",X"7F",X"DD",X"DA",X"FF",
		X"7F",X"DD",X"DA",X"FF",X"7F",X"DD",X"DA",X"FF",X"7F",X"DD",X"DA",X"FF",X"7F",X"DD",X"DA",X"FF",
		X"7F",X"DD",X"DA",X"FF",X"7F",X"DD",X"DA",X"FF",X"7F",X"DD",X"DA",X"FF",X"7F",X"DD",X"DA",X"FF",
		X"7F",X"DD",X"DA",X"FF",X"7F",X"DD",X"DA",X"FF",X"7F",X"DD",X"DA",X"FF",X"7F",X"DD",X"DA",X"FF",
		X"99",X"99",X"99",X"99",X"FF",X"FF",X"FF",X"FF",X"75",X"F5",X"FF",X"5F",X"7F",X"F5",X"FF",X"5F",
		X"7F",X"F5",X"FF",X"5F",X"FF",X"F5",X"FF",X"5F",X"5F",X"55",X"55",X"55",X"5F",X"55",X"55",X"55",
		X"FF",X"F2",X"FF",X"FF",X"FF",X"5F",X"2F",X"7F",X"5F",X"55",X"F5",X"7F",X"5F",X"55",X"55",X"F5",
		X"5F",X"55",X"5F",X"5F",X"5F",X"55",X"FF",X"F5",X"5F",X"55",X"2F",X"FF",X"FF",X"55",X"2F",X"77",
		X"77",X"AA",X"22",X"F7",X"77",X"AA",X"22",X"F7",X"77",X"FF",X"CC",X"F7",X"EE",X"FF",X"CC",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"CF",X"FF",X"FF",X"FC",X"7F",X"AA",X"FF",X"FF",X"7F",X"EE",X"FF",X"AF",
		X"7F",X"77",X"C7",X"77",X"7F",X"77",X"77",X"77",X"7F",X"FF",X"FF",X"77",X"7F",X"AA",X"AA",X"77",
		X"7F",X"CC",X"CC",X"7F",X"FF",X"CC",X"CC",X"77",X"CF",X"CC",X"CC",X"8F",X"7F",X"22",X"22",X"FC");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
