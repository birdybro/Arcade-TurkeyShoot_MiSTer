library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity turkey_shoot_sound is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of turkey_shoot_sound is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"EA",X"0F",X"8E",X"00",X"FF",X"CE",X"20",X"00",X"6F",X"01",X"6F",X"03",X"86",X"FF",X"A7",X"02",
		X"6F",X"00",X"86",X"37",X"A7",X"01",X"86",X"3C",X"A7",X"03",X"CE",X"00",X"FF",X"6F",X"00",X"09",
		X"26",X"FB",X"7A",X"00",X"81",X"7A",X"00",X"80",X"7A",X"00",X"80",X"0E",X"20",X"09",X"8E",X"00",
		X"FF",X"B6",X"20",X"00",X"0E",X"8D",X"28",X"86",X"3C",X"B7",X"20",X"03",X"86",X"37",X"B7",X"20",
		X"01",X"20",X"FE",X"0F",X"8E",X"00",X"FF",X"4F",X"CE",X"FF",X"FF",X"5F",X"E9",X"00",X"09",X"8C",
		X"E0",X"00",X"26",X"F8",X"E1",X"00",X"26",X"FE",X"86",X"55",X"8D",X"03",X"20",X"FA",X"39",X"C6",
		X"3C",X"F7",X"20",X"03",X"C6",X"3F",X"F7",X"20",X"01",X"81",X"01",X"25",X"F1",X"81",X"18",X"22",
		X"07",X"4A",X"BD",X"E0",X"E0",X"7E",X"E1",X"46",X"81",X"2F",X"22",X"05",X"80",X"19",X"7E",X"F2",
		X"BD",X"81",X"4E",X"22",X"0D",X"80",X"30",X"CE",X"E0",X"A2",X"48",X"BD",X"F1",X"1A",X"EE",X"00",
		X"6E",X"00",X"81",X"56",X"22",X"05",X"80",X"4F",X"7E",X"EF",X"87",X"81",X"57",X"22",X"BF",X"7E",
		X"FB",X"4B",X"E4",X"FE",X"E5",X"09",X"E5",X"A3",X"E6",X"65",X"E5",X"1C",X"E5",X"20",X"E5",X"24",
		X"E6",X"6D",X"E6",X"75",X"E6",X"F4",X"E7",X"8E",X"E7",X"F9",X"E8",X"0B",X"E8",X"9E",X"F4",X"D6",
		X"F1",X"29",X"E8",X"D3",X"E8",X"D7",X"E8",X"DB",X"E8",X"DF",X"F1",X"41",X"F1",X"65",X"F1",X"8F",
		X"F1",X"9E",X"F1",X"B7",X"F1",X"F0",X"F2",X"0F",X"F2",X"60",X"F2",X"C2",X"E7",X"6B",X"F2",X"A4",
		X"16",X"58",X"1B",X"1B",X"1B",X"CE",X"E3",X"5D",X"BD",X"F1",X"1A",X"A6",X"00",X"16",X"84",X"0F",
		X"97",X"95",X"54",X"54",X"54",X"54",X"D7",X"94",X"A6",X"01",X"16",X"54",X"54",X"54",X"54",X"D7",
		X"96",X"84",X"0F",X"97",X"87",X"DF",X"8A",X"CE",X"E2",X"25",X"7A",X"00",X"87",X"2B",X"08",X"A6",
		X"00",X"4C",X"BD",X"F1",X"1A",X"20",X"F3",X"DF",X"99",X"BD",X"E1",X"D0",X"DE",X"8A",X"A6",X"02",
		X"97",X"9B",X"BD",X"E1",X"E2",X"DE",X"8A",X"A6",X"03",X"97",X"97",X"A6",X"04",X"97",X"98",X"A6",
		X"05",X"16",X"A6",X"06",X"CE",X"E4",X"0C",X"BD",X"F1",X"1A",X"17",X"DF",X"9C",X"7F",X"00",X"A4",
		X"BD",X"F1",X"1A",X"DF",X"9E",X"39",X"96",X"94",X"97",X"A3",X"DE",X"9C",X"DF",X"8C",X"DE",X"8C",
		X"A6",X"00",X"9B",X"A4",X"97",X"A2",X"9C",X"9E",X"27",X"26",X"D6",X"95",X"08",X"DF",X"8C",X"CE",
		X"00",X"A5",X"96",X"A2",X"4A",X"26",X"FD",X"A6",X"00",X"B7",X"20",X"02",X"08",X"9C",X"A0",X"26",
		X"F1",X"5A",X"27",X"DA",X"08",X"09",X"08",X"09",X"08",X"09",X"08",X"09",X"01",X"01",X"20",X"DF",
		X"96",X"96",X"8D",X"5E",X"7A",X"00",X"A3",X"26",X"C1",X"96",X"97",X"27",X"42",X"7A",X"00",X"98",
		X"27",X"3D",X"9B",X"A4",X"97",X"A4",X"DE",X"9C",X"5F",X"96",X"A4",X"7D",X"00",X"97",X"2B",X"06",
		X"AB",X"00",X"25",X"08",X"20",X"0B",X"AB",X"00",X"27",X"02",X"25",X"05",X"5D",X"27",X"08",X"20",
		X"0F",X"5D",X"26",X"03",X"DF",X"9C",X"5C",X"08",X"9C",X"9E",X"26",X"DD",X"5D",X"26",X"01",X"39",
		X"DF",X"9E",X"96",X"96",X"27",X"06",X"8D",X"08",X"96",X"9B",X"8D",X"16",X"7E",X"E1",X"46",X"39",
		X"CE",X"00",X"A5",X"DF",X"8E",X"DE",X"99",X"E6",X"00",X"08",X"BD",X"E2",X"11",X"DE",X"8E",X"DF",
		X"A0",X"39",X"4D",X"27",X"2B",X"DE",X"99",X"DF",X"8C",X"CE",X"00",X"A5",X"97",X"88",X"DF",X"8E",
		X"DE",X"8C",X"D6",X"88",X"D7",X"87",X"E6",X"01",X"54",X"54",X"54",X"54",X"08",X"DF",X"8C",X"DE",
		X"8E",X"A6",X"00",X"10",X"7A",X"00",X"87",X"26",X"FA",X"A7",X"00",X"08",X"9C",X"A0",X"26",X"DE",
		X"39",X"36",X"A6",X"00",X"DF",X"8C",X"DE",X"8E",X"A7",X"00",X"08",X"DF",X"8E",X"DE",X"8C",X"08",
		X"5A",X"26",X"EF",X"32",X"39",X"08",X"7F",X"D9",X"FF",X"D9",X"7F",X"24",X"00",X"24",X"08",X"00",
		X"40",X"80",X"00",X"FF",X"00",X"80",X"40",X"10",X"7F",X"B0",X"D9",X"F5",X"FF",X"F5",X"D9",X"B0",
		X"7F",X"4E",X"24",X"09",X"00",X"09",X"24",X"4E",X"10",X"7F",X"C5",X"EC",X"E7",X"BF",X"8D",X"6D",
		X"6A",X"7F",X"94",X"92",X"71",X"40",X"17",X"12",X"39",X"10",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"48",X"8A",X"95",X"A0",X"AB",X"B5",
		X"BF",X"C8",X"D1",X"DA",X"E1",X"E8",X"EE",X"F3",X"F7",X"FB",X"FD",X"FE",X"FF",X"FE",X"FD",X"FB",
		X"F7",X"F3",X"EE",X"E8",X"E1",X"DA",X"D1",X"C8",X"BF",X"B5",X"AB",X"A0",X"95",X"8A",X"7F",X"75",
		X"6A",X"5F",X"54",X"4A",X"40",X"37",X"2E",X"25",X"1E",X"17",X"11",X"0C",X"08",X"04",X"02",X"01",
		X"00",X"01",X"02",X"04",X"08",X"0C",X"11",X"17",X"1E",X"25",X"2E",X"37",X"40",X"4A",X"54",X"5F",
		X"6A",X"75",X"7F",X"10",X"59",X"7B",X"98",X"AC",X"B3",X"AC",X"98",X"7B",X"59",X"37",X"19",X"06",
		X"00",X"06",X"19",X"37",X"08",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"10",X"76",X"FF",
		X"B8",X"D0",X"9D",X"E6",X"6A",X"82",X"76",X"EA",X"81",X"86",X"4E",X"9C",X"32",X"63",X"10",X"00",
		X"F4",X"00",X"E8",X"00",X"DC",X"00",X"E2",X"00",X"DC",X"00",X"E8",X"00",X"F4",X"00",X"00",X"1C",
		X"80",X"40",X"29",X"1B",X"10",X"09",X"06",X"04",X"07",X"0C",X"12",X"1E",X"30",X"49",X"A4",X"C9",
		X"DF",X"EB",X"F6",X"FB",X"FF",X"FF",X"FB",X"F5",X"EA",X"DD",X"C7",X"9B",X"0C",X"00",X"50",X"60",
		X"B0",X"20",X"20",X"F0",X"90",X"80",X"C0",X"50",X"70",X"10",X"3C",X"10",X"17",X"3F",X"70",X"92",
		X"95",X"7F",X"7C",X"7E",X"8A",X"BE",X"E7",X"EF",X"C5",X"7F",X"08",X"00",X"20",X"40",X"60",X"80",
		X"A0",X"C0",X"E0",X"08",X"FF",X"DF",X"BF",X"9F",X"7F",X"5F",X"3F",X"1F",X"20",X"4C",X"45",X"41",
		X"41",X"43",X"47",X"77",X"87",X"90",X"97",X"A1",X"A7",X"AE",X"B5",X"B8",X"BC",X"BE",X"BF",X"C1",
		X"C2",X"C2",X"C2",X"C1",X"BF",X"BE",X"BB",X"B6",X"B1",X"AC",X"A4",X"9E",X"93",X"F6",X"57",X"00",
		X"00",X"02",X"06",X"9E",X"73",X"2A",X"00",X"00",X"00",X"04",X"08",X"14",X"0A",X"00",X"00",X"00",
		X"04",X"00",X"14",X"0A",X"00",X"00",X"00",X"04",X"04",X"14",X"02",X"00",X"00",X"00",X"09",X"0C",
		X"11",X"02",X"00",X"00",X"00",X"28",X"15",X"1F",X"0B",X"00",X"00",X"00",X"0F",X"3D",X"18",X"00",
		X"00",X"02",X"01",X"20",X"4C",X"11",X"02",X"00",X"00",X"00",X"18",X"6C",X"15",X"02",X"00",X"00",
		X"00",X"16",X"84",X"81",X"02",X"00",X"00",X"00",X"04",X"9A",X"11",X"12",X"00",X"00",X"00",X"63",
		X"00",X"11",X"15",X"00",X"00",X"00",X"63",X"00",X"11",X"10",X"00",X"00",X"00",X"63",X"00",X"11",
		X"11",X"00",X"00",X"00",X"63",X"00",X"16",X"02",X"00",X"00",X"00",X"7C",X"3D",X"1F",X"0C",X"00",
		X"FF",X"30",X"09",X"0C",X"F1",X"19",X"00",X"00",X"00",X"20",X"43",X"52",X"36",X"00",X"00",X"00",
		X"10",X"BB",X"A3",X"19",X"00",X"01",X"01",X"10",X"CB",X"16",X"82",X"00",X"0E",X"01",X"0E",X"DB",
		X"63",X"26",X"00",X"00",X"00",X"10",X"CB",X"23",X"15",X"00",X"02",X"07",X"03",X"E9",X"82",X"19",
		X"00",X"01",X"01",X"20",X"43",X"82",X"15",X"00",X"03",X"01",X"20",X"43",X"20",X"18",X"20",X"01",
		X"01",X"30",X"28",X"30",X"08",X"10",X"20",X"30",X"20",X"10",X"0C",X"0A",X"08",X"07",X"06",X"05",
		X"04",X"60",X"45",X"28",X"21",X"5D",X"42",X"25",X"1E",X"58",X"3D",X"20",X"19",X"60",X"38",X"28",
		X"14",X"4C",X"31",X"14",X"0D",X"40",X"25",X"08",X"01",X"4C",X"31",X"14",X"0D",X"40",X"25",X"08",
		X"01",X"4C",X"31",X"14",X"0D",X"40",X"25",X"08",X"01",X"0A",X"09",X"08",X"07",X"06",X"05",X"06",
		X"07",X"08",X"09",X"0A",X"0A",X"0A",X"0A",X"0A",X"20",X"1F",X"1E",X"1D",X"1C",X"1B",X"1A",X"19",
		X"18",X"17",X"16",X"15",X"14",X"13",X"12",X"11",X"10",X"0F",X"0E",X"0D",X"0C",X"0B",X"0A",X"09",
		X"08",X"07",X"06",X"05",X"05",X"05",X"05",X"05",X"60",X"45",X"28",X"21",X"58",X"3D",X"20",X"19",
		X"4C",X"31",X"14",X"0D",X"40",X"25",X"08",X"01",X"34",X"1C",X"08",X"01",X"28",X"15",X"08",X"01",
		X"1E",X"02",X"1B",X"04",X"23",X"07",X"1D",X"01",X"22",X"03",X"19",X"09",X"1F",X"06",X"1A",X"05",
		X"1C",X"0B",X"21",X"08",X"20",X"0A",X"60",X"45",X"28",X"21",X"07",X"08",X"09",X"0A",X"0C",X"08",
		X"01",X"40",X"02",X"42",X"03",X"43",X"04",X"44",X"05",X"45",X"06",X"46",X"07",X"47",X"08",X"48",
		X"09",X"49",X"0A",X"4A",X"0B",X"4B",X"00",X"01",X"01",X"02",X"02",X"04",X"04",X"08",X"08",X"10",
		X"20",X"28",X"30",X"38",X"40",X"48",X"50",X"14",X"18",X"20",X"30",X"40",X"50",X"40",X"30",X"20",
		X"10",X"0C",X"0A",X"08",X"07",X"06",X"05",X"0C",X"08",X"80",X"10",X"78",X"18",X"70",X"20",X"60",
		X"28",X"58",X"30",X"50",X"40",X"10",X"08",X"01",X"01",X"01",X"01",X"FF",X"03",X"E8",X"CE",X"E4",
		X"F8",X"20",X"09",X"01",X"01",X"01",X"40",X"10",X"00",X"CE",X"E5",X"03",X"A6",X"00",X"97",X"99",
		X"A6",X"01",X"97",X"9A",X"A6",X"02",X"E6",X"03",X"EE",X"04",X"20",X"0F",X"C6",X"02",X"20",X"06",
		X"C6",X"03",X"20",X"02",X"C6",X"04",X"4F",X"97",X"9A",X"97",X"99",X"97",X"98",X"D7",X"93",X"DF",
		X"96",X"7F",X"00",X"95",X"DE",X"96",X"B6",X"20",X"02",X"16",X"54",X"54",X"54",X"D8",X"81",X"54",
		X"76",X"00",X"80",X"76",X"00",X"81",X"D6",X"93",X"7D",X"00",X"99",X"27",X"04",X"D4",X"80",X"DB",
		X"9A",X"D7",X"94",X"D6",X"95",X"91",X"81",X"22",X"12",X"09",X"27",X"26",X"B7",X"20",X"02",X"DB",
		X"95",X"99",X"94",X"25",X"16",X"91",X"81",X"23",X"F0",X"20",X"10",X"09",X"27",X"14",X"B7",X"20",
		X"02",X"D0",X"95",X"92",X"94",X"25",X"04",X"91",X"81",X"22",X"F0",X"96",X"81",X"B7",X"20",X"02",
		X"20",X"B7",X"D6",X"98",X"27",X"B3",X"96",X"93",X"D6",X"95",X"44",X"56",X"44",X"56",X"44",X"56",
		X"43",X"50",X"82",X"FF",X"DB",X"95",X"99",X"93",X"D7",X"95",X"97",X"93",X"26",X"96",X"C1",X"07",
		X"26",X"92",X"39",X"7F",X"20",X"02",X"CE",X"10",X"00",X"09",X"26",X"FD",X"39",X"CE",X"E6",X"61",
		X"DF",X"84",X"CE",X"00",X"93",X"DF",X"8E",X"C6",X"AF",X"D7",X"89",X"39",X"DF",X"8C",X"CE",X"E6",
		X"61",X"DF",X"84",X"86",X"80",X"D6",X"96",X"2A",X"09",X"D6",X"81",X"54",X"54",X"54",X"5C",X"5A",
		X"26",X"FD",X"7A",X"00",X"9B",X"27",X"4C",X"7A",X"00",X"9C",X"27",X"4C",X"7A",X"00",X"9D",X"27",
		X"4C",X"7A",X"00",X"9E",X"26",X"DF",X"D6",X"96",X"27",X"DB",X"C4",X"7F",X"D7",X"9E",X"D6",X"81",
		X"58",X"DB",X"81",X"CB",X"0B",X"D7",X"81",X"7A",X"00",X"AE",X"26",X"0E",X"D6",X"A2",X"D7",X"AE",
		X"DE",X"84",X"09",X"8C",X"E6",X"5A",X"27",X"4E",X"DF",X"84",X"D6",X"81",X"2B",X"06",X"D4",X"9A",
		X"C4",X"7F",X"20",X"05",X"D4",X"9A",X"C4",X"7F",X"50",X"36",X"1B",X"16",X"32",X"DE",X"84",X"AD",
		X"00",X"20",X"A2",X"CE",X"00",X"93",X"20",X"08",X"CE",X"00",X"94",X"20",X"03",X"CE",X"00",X"95",
		X"6D",X"18",X"27",X"12",X"6A",X"18",X"26",X"0E",X"E6",X"0C",X"E7",X"18",X"E6",X"00",X"EB",X"10",
		X"E1",X"14",X"27",X"12",X"E7",X"00",X"E6",X"00",X"E7",X"08",X"AB",X"04",X"60",X"04",X"16",X"DE",
		X"84",X"AD",X"00",X"7E",X"E5",X"C5",X"DE",X"8C",X"39",X"54",X"54",X"54",X"54",X"54",X"54",X"54",
		X"54",X"F7",X"20",X"02",X"39",X"BD",X"E5",X"AD",X"CE",X"E6",X"D8",X"20",X"0E",X"BD",X"E5",X"AD",
		X"CE",X"E6",X"BC",X"20",X"06",X"BD",X"E5",X"AD",X"CE",X"E6",X"A0",X"C6",X"1C",X"BD",X"E2",X"11",
		X"7E",X"E5",X"BC",X"39",X"FF",X"FF",X"FF",X"90",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"90",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"00",X"00",X"00",X"7F",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"7F",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"04",X"00",X"00",X"04",
		X"7F",X"00",X"00",X"7F",X"04",X"00",X"00",X"04",X"FF",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"A0",X"02",X"80",X"00",X"30",X"0A",X"7F",X"00",X"7F",
		X"02",X"80",X"00",X"30",X"C0",X"80",X"00",X"20",X"01",X"10",X"00",X"15",X"C0",X"10",X"00",X"00",
		X"C0",X"80",X"00",X"00",X"BD",X"E5",X"AD",X"86",X"80",X"97",X"9D",X"86",X"E7",X"97",X"9B",X"86",
		X"80",X"97",X"87",X"86",X"12",X"4A",X"26",X"FD",X"96",X"9A",X"9B",X"9D",X"97",X"9A",X"44",X"44",
		X"44",X"8B",X"2B",X"97",X"9C",X"DE",X"9B",X"A6",X"00",X"B7",X"20",X"02",X"7A",X"00",X"87",X"26",
		X"E2",X"7A",X"00",X"9D",X"96",X"9D",X"81",X"20",X"26",X"D5",X"39",X"80",X"8C",X"98",X"A5",X"B0",
		X"BC",X"C6",X"D0",X"DA",X"E2",X"EA",X"F0",X"F5",X"FA",X"FD",X"FE",X"FF",X"FE",X"FD",X"FA",X"F5",
		X"F0",X"EA",X"E2",X"DA",X"D0",X"C6",X"BC",X"B0",X"A5",X"98",X"8C",X"80",X"73",X"67",X"5A",X"4F",
		X"43",X"39",X"2F",X"25",X"1D",X"15",X"0F",X"0A",X"05",X"02",X"01",X"00",X"01",X"02",X"05",X"0A",
		X"0F",X"15",X"1D",X"25",X"2F",X"39",X"43",X"4F",X"5A",X"67",X"73",X"86",X"30",X"B7",X"20",X"02",
		X"CE",X"01",X"20",X"86",X"48",X"4A",X"26",X"FD",X"73",X"20",X"02",X"09",X"26",X"F5",X"CE",X"01",
		X"20",X"86",X"58",X"4A",X"26",X"FD",X"73",X"20",X"02",X"09",X"26",X"F5",X"20",X"E2",X"7F",X"20",
		X"04",X"CE",X"E7",X"D5",X"DF",X"95",X"DE",X"95",X"A6",X"00",X"27",X"33",X"E6",X"01",X"C4",X"F0",
		X"D7",X"94",X"E6",X"01",X"08",X"08",X"DF",X"95",X"97",X"93",X"C4",X"0F",X"96",X"94",X"B7",X"20",
		X"02",X"96",X"93",X"CE",X"00",X"05",X"09",X"26",X"FD",X"4A",X"26",X"F7",X"7F",X"20",X"02",X"96",
		X"93",X"CE",X"00",X"05",X"09",X"26",X"FD",X"4A",X"26",X"F7",X"5A",X"26",X"DF",X"20",X"C7",X"86",
		X"80",X"B7",X"20",X"04",X"39",X"01",X"FC",X"02",X"FC",X"03",X"F8",X"04",X"F8",X"06",X"F8",X"08",
		X"F4",X"0C",X"F4",X"10",X"F4",X"20",X"F2",X"40",X"F1",X"60",X"F1",X"80",X"F1",X"A0",X"F1",X"C0",
		X"F1",X"00",X"00",X"FE",X"04",X"02",X"04",X"FF",X"00",X"BD",X"E5",X"AD",X"CE",X"E7",X"F3",X"BD",
		X"E8",X"2A",X"7E",X"E8",X"43",X"50",X"FF",X"00",X"00",X"60",X"80",X"BD",X"E5",X"AD",X"C6",X"30",
		X"CE",X"E8",X"05",X"8D",X"15",X"96",X"81",X"48",X"9B",X"81",X"8B",X"0B",X"97",X"81",X"44",X"44",
		X"8B",X"0C",X"97",X"94",X"8D",X"1D",X"5A",X"26",X"EC",X"39",X"A6",X"00",X"97",X"94",X"A6",X"01",
		X"97",X"95",X"A6",X"02",X"97",X"96",X"A6",X"03",X"97",X"97",X"A6",X"04",X"97",X"98",X"A6",X"05",
		X"97",X"99",X"39",X"96",X"89",X"37",X"D6",X"98",X"D7",X"9A",X"D6",X"95",X"D7",X"9B",X"43",X"D6",
		X"94",X"B7",X"20",X"02",X"5A",X"26",X"FD",X"43",X"D6",X"94",X"20",X"00",X"08",X"09",X"08",X"09",
		X"B7",X"20",X"02",X"5A",X"26",X"FD",X"7A",X"00",X"9B",X"27",X"16",X"7A",X"00",X"9A",X"26",X"DE",
		X"43",X"D6",X"98",X"B7",X"20",X"02",X"D7",X"9A",X"D6",X"94",X"9B",X"99",X"2B",X"1E",X"01",X"20",
		X"15",X"08",X"09",X"01",X"43",X"D6",X"95",X"B7",X"20",X"02",X"D7",X"9B",X"D6",X"94",X"D0",X"96",
		X"D1",X"97",X"D1",X"97",X"27",X"06",X"D7",X"94",X"C0",X"05",X"20",X"B8",X"33",X"39",X"86",X"01",
		X"97",X"9A",X"C6",X"03",X"97",X"99",X"86",X"FF",X"B7",X"20",X"02",X"D7",X"95",X"D6",X"95",X"96",
		X"81",X"44",X"44",X"44",X"98",X"81",X"44",X"76",X"00",X"80",X"76",X"00",X"81",X"24",X"03",X"73",
		X"20",X"02",X"96",X"99",X"4A",X"26",X"FD",X"5A",X"26",X"E5",X"96",X"99",X"9B",X"9A",X"97",X"99",
		X"26",X"DB",X"39",X"86",X"00",X"20",X"29",X"86",X"01",X"20",X"25",X"86",X"02",X"20",X"21",X"86",
		X"03",X"8D",X"1D",X"86",X"04",X"20",X"19",X"0D",X"40",X"F0",X"FF",X"12",X"08",X"A8",X"18",X"01",
		X"08",X"04",X"A8",X"18",X"01",X"10",X"04",X"20",X"F8",X"FF",X"20",X"10",X"F0",X"10",X"01",X"01",
		X"CE",X"D9",X"39",X"DF",X"80",X"16",X"48",X"48",X"1B",X"CE",X"E8",X"E7",X"BD",X"F1",X"1A",X"A6",
		X"00",X"97",X"AB",X"A6",X"01",X"97",X"94",X"A6",X"02",X"97",X"93",X"A6",X"03",X"97",X"98",X"A6",
		X"04",X"97",X"B0",X"8D",X"30",X"8D",X"58",X"96",X"AF",X"91",X"B0",X"26",X"F8",X"59",X"F7",X"20",
		X"02",X"8D",X"2D",X"8D",X"38",X"8D",X"5C",X"7D",X"00",X"94",X"27",X"23",X"7D",X"00",X"95",X"26",
		X"E4",X"7D",X"00",X"98",X"27",X"DF",X"2B",X"05",X"7C",X"00",X"B0",X"20",X"D8",X"7A",X"00",X"B0",
		X"7A",X"00",X"AF",X"20",X"D0",X"7F",X"00",X"95",X"96",X"B0",X"97",X"AF",X"7F",X"00",X"AE",X"39",
		X"96",X"81",X"44",X"44",X"44",X"98",X"81",X"97",X"A9",X"08",X"84",X"07",X"39",X"96",X"A9",X"44",
		X"76",X"00",X"80",X"76",X"00",X"81",X"86",X"00",X"24",X"02",X"96",X"94",X"97",X"AE",X"39",X"96",
		X"B0",X"7A",X"00",X"AF",X"27",X"04",X"08",X"09",X"20",X"08",X"97",X"AF",X"D6",X"AE",X"54",X"7C",
		X"00",X"95",X"39",X"96",X"AB",X"91",X"95",X"27",X"04",X"08",X"09",X"20",X"09",X"7F",X"00",X"95",
		X"96",X"94",X"90",X"93",X"97",X"94",X"39",X"C0",X"0D",X"37",X"BD",X"00",X"AC",X"33",X"C1",X"14",
		X"22",X"F5",X"01",X"96",X"A4",X"9B",X"A1",X"97",X"A4",X"C9",X"F6",X"5A",X"2A",X"FD",X"96",X"A8",
		X"4C",X"84",X"0F",X"8A",X"90",X"97",X"A8",X"DE",X"A7",X"E6",X"00",X"F7",X"20",X"02",X"84",X"0F",
		X"39",X"4F",X"CE",X"00",X"90",X"C6",X"61",X"A7",X"00",X"08",X"5A",X"26",X"FA",X"C6",X"DF",X"D7",
		X"A6",X"C6",X"B7",X"D7",X"B0",X"C6",X"7E",X"D7",X"AC",X"CE",X"EB",X"BC",X"DF",X"AD",X"D6",X"8C",
		X"D7",X"A3",X"C0",X"03",X"BD",X"E9",X"AE",X"08",X"D6",X"A3",X"C0",X"02",X"BD",X"E9",X"A7",X"26",
		X"F7",X"D6",X"A0",X"96",X"A1",X"9B",X"8D",X"D9",X"8C",X"97",X"8D",X"D7",X"8C",X"DB",X"A2",X"86",
		X"19",X"11",X"24",X"01",X"81",X"16",X"D7",X"A3",X"01",X"C0",X"09",X"BD",X"E9",X"AE",X"96",X"AF",
		X"16",X"48",X"C9",X"00",X"D7",X"AF",X"D6",X"A3",X"C0",X"05",X"96",X"A5",X"2A",X"06",X"7C",X"00",
		X"A5",X"01",X"20",X"BE",X"5A",X"BD",X"E9",X"AE",X"DE",X"8A",X"A6",X"00",X"2A",X"12",X"81",X"80",
		X"27",X"5F",X"4C",X"97",X"A5",X"08",X"FF",X"00",X"8A",X"D6",X"A3",X"C0",X"06",X"7E",X"E9",X"F2",
		X"08",X"E6",X"00",X"37",X"08",X"DF",X"8A",X"97",X"A9",X"84",X"70",X"44",X"44",X"44",X"5F",X"8B",
		X"35",X"C9",X"EB",X"97",X"AB",X"D7",X"AA",X"D6",X"A3",X"D6",X"A3",X"C0",X"0D",X"BD",X"E9",X"AE",
		X"5F",X"DE",X"AA",X"EE",X"00",X"6E",X"00",X"96",X"A9",X"47",X"C2",X"00",X"D4",X"8C",X"32",X"10",
		X"9B",X"8C",X"97",X"8C",X"08",X"D6",X"A3",X"C0",X"0A",X"7E",X"E9",X"F4",X"96",X"A9",X"47",X"C2",
		X"00",X"D4",X"A2",X"32",X"10",X"9B",X"A2",X"97",X"A2",X"20",X"EA",X"32",X"DE",X"8A",X"09",X"6E",
		X"00",X"96",X"A6",X"81",X"DF",X"2B",X"01",X"39",X"D6",X"A3",X"C0",X"07",X"BD",X"E9",X"AE",X"DE",
		X"A5",X"6A",X"02",X"2B",X"12",X"EE",X"00",X"A6",X"00",X"36",X"08",X"DF",X"8A",X"F6",X"00",X"A3",
		X"C0",X"09",X"BD",X"E9",X"AE",X"20",X"55",X"EE",X"00",X"08",X"DF",X"8A",X"96",X"A6",X"8B",X"03",
		X"97",X"A6",X"D6",X"A3",X"C0",X"07",X"01",X"7E",X"E9",X"F2",X"08",X"20",X"04",X"D7",X"A0",X"D7",
		X"A1",X"D6",X"A9",X"C4",X"0F",X"CB",X"F8",X"C8",X"F8",X"32",X"9B",X"A1",X"D9",X"A0",X"97",X"A1",
		X"D7",X"A0",X"F6",X"00",X"A3",X"C0",X"09",X"7E",X"E9",X"F2",X"96",X"A6",X"80",X"03",X"97",X"A6",
		X"DE",X"A5",X"96",X"8B",X"D6",X"8A",X"8B",X"FF",X"C9",X"FF",X"E7",X"00",X"A7",X"01",X"D6",X"A9",
		X"C4",X"0F",X"E7",X"02",X"D6",X"A3",X"C0",X"0C",X"BD",X"E9",X"AE",X"08",X"08",X"08",X"5F",X"01",
		X"32",X"47",X"49",X"C2",X"00",X"9B",X"8B",X"D9",X"8A",X"97",X"8B",X"F7",X"00",X"8A",X"D6",X"A3",
		X"C0",X"07",X"7E",X"E9",X"F2",X"EA",X"77",X"EA",X"8C",X"EA",X"DD",X"EA",X"DA",X"EA",X"77",X"EA",
		X"9B",X"EA",X"FA",X"EB",X"20",X"EC",X"B9",X"ED",X"42",X"EB",X"F1",X"EC",X"EA",X"EB",X"6C",X"EC",
		X"FB",X"EB",X"97",X"EC",X"2E",X"DE",X"AF",X"EE",X"03",X"08",X"DF",X"88",X"BD",X"EC",X"28",X"08",
		X"39",X"EE",X"00",X"DF",X"88",X"CE",X"EC",X"2E",X"DF",X"AD",X"01",X"39",X"96",X"B0",X"81",X"B7",
		X"23",X"12",X"DE",X"AF",X"6A",X"02",X"2A",X"E9",X"80",X"03",X"97",X"B0",X"CE",X"EB",X"55",X"DF",
		X"AD",X"6D",X"00",X"39",X"CE",X"EB",X"8C",X"DF",X"AD",X"01",X"20",X"05",X"08",X"08",X"01",X"8D",
		X"05",X"8D",X"03",X"6D",X"00",X"01",X"39",X"DE",X"AF",X"96",X"88",X"A7",X"03",X"96",X"89",X"A7",
		X"04",X"96",X"B9",X"84",X"0F",X"A7",X"05",X"08",X"CE",X"EB",X"AE",X"DF",X"AD",X"39",X"96",X"B0",
		X"8B",X"03",X"97",X"B0",X"CE",X"EC",X"2E",X"DF",X"AD",X"01",X"20",X"D5",X"7D",X"00",X"AF",X"26",
		X"CE",X"DE",X"88",X"A6",X"00",X"08",X"DF",X"88",X"97",X"B9",X"2A",X"05",X"97",X"AF",X"A6",X"00",
		X"39",X"CE",X"EB",X"D8",X"FF",X"00",X"AD",X"39",X"5F",X"96",X"B9",X"84",X"70",X"44",X"44",X"44",
		X"8B",X"45",X"C9",X"EB",X"D7",X"B7",X"97",X"B8",X"DE",X"B7",X"EE",X"00",X"DF",X"AD",X"DF",X"AD",
		X"39",X"96",X"B9",X"84",X"0F",X"4C",X"4C",X"97",X"AF",X"20",X"1D",X"7C",X"00",X"B2",X"DE",X"B1",
		X"8C",X"00",X"E8",X"27",X"13",X"A6",X"00",X"CE",X"EC",X"42",X"97",X"B5",X"27",X"03",X"7E",X"EC",
		X"14",X"CE",X"EB",X"FB",X"DF",X"AD",X"08",X"39",X"86",X"DE",X"B7",X"00",X"B2",X"CE",X"EB",X"FB",
		X"7A",X"00",X"AF",X"27",X"03",X"7E",X"EC",X"2B",X"CE",X"EB",X"BC",X"DF",X"AD",X"39",X"DE",X"88",
		X"5F",X"A6",X"00",X"4C",X"47",X"49",X"C2",X"00",X"9B",X"89",X"D9",X"88",X"97",X"89",X"D7",X"88",
		X"20",X"E6",X"96",X"B2",X"80",X"DF",X"48",X"5F",X"9B",X"8F",X"D9",X"8E",X"D7",X"B7",X"97",X"B8",
		X"86",X"80",X"97",X"B6",X"CE",X"EC",X"5F",X"DF",X"AD",X"CE",X"00",X"90",X"DF",X"B3",X"39",X"DE",
		X"B7",X"EE",X"00",X"DF",X"B7",X"CE",X"EC",X"74",X"DF",X"AD",X"DE",X"B1",X"A6",X"09",X"9B",X"B5",
		X"A7",X"09",X"08",X"39",X"96",X"B6",X"27",X"1D",X"74",X"00",X"B6",X"DE",X"B3",X"E6",X"00",X"94",
		X"B7",X"26",X"09",X"FB",X"00",X"B5",X"E7",X"00",X"7C",X"00",X"B4",X"39",X"F0",X"00",X"B5",X"E7",
		X"00",X"7C",X"00",X"B4",X"39",X"D6",X"B4",X"C1",X"A0",X"27",X"0B",X"D6",X"B8",X"D7",X"B7",X"C6",
		X"80",X"F7",X"00",X"B6",X"20",X"0F",X"CE",X"EB",X"BC",X"D6",X"AF",X"26",X"03",X"7E",X"EC",X"B3",
		X"CE",X"EB",X"FB",X"DF",X"AD",X"6D",X"00",X"08",X"39",X"96",X"B9",X"84",X"07",X"8B",X"E0",X"97",
		X"B2",X"DE",X"88",X"A6",X"00",X"08",X"DF",X"88",X"97",X"B5",X"CE",X"EC",X"D1",X"DF",X"AD",X"08",
		X"39",X"DE",X"B1",X"5F",X"96",X"B9",X"8B",X"F8",X"C2",X"00",X"E4",X"09",X"50",X"DB",X"B5",X"D7",
		X"B5",X"CE",X"EC",X"42",X"DF",X"AD",X"08",X"08",X"01",X"39",X"D6",X"B9",X"54",X"C4",X"07",X"CA",
		X"E0",X"D7",X"B2",X"C6",X"FF",X"C9",X"00",X"C9",X"00",X"20",X"E4",X"96",X"B9",X"47",X"25",X"13",
		X"CE",X"00",X"00",X"DF",X"E0",X"DF",X"E2",X"DF",X"E4",X"DF",X"E6",X"08",X"CE",X"EB",X"BC",X"FF",
		X"00",X"AD",X"39",X"85",X"02",X"26",X"0C",X"C6",X"DF",X"D7",X"B2",X"CE",X"ED",X"28",X"DF",X"AD",
		X"7E",X"EB",X"93",X"FE",X"00",X"88",X"20",X"F6",X"5F",X"96",X"B9",X"8B",X"AE",X"C2",X"00",X"D4",
		X"E8",X"DE",X"88",X"A6",X"00",X"08",X"DF",X"88",X"10",X"97",X"B5",X"CE",X"EC",X"42",X"FF",X"00",
		X"AD",X"39",X"C6",X"E0",X"D7",X"B2",X"DE",X"88",X"E6",X"00",X"D7",X"B7",X"08",X"DF",X"88",X"D6",
		X"B9",X"54",X"24",X"18",X"CE",X"ED",X"86",X"DF",X"AD",X"39",X"5F",X"96",X"B8",X"47",X"C2",X"00",
		X"DE",X"B1",X"E4",X"00",X"1B",X"A7",X"00",X"7C",X"00",X"B2",X"A6",X"00",X"CE",X"ED",X"72",X"DF",
		X"AD",X"39",X"78",X"00",X"B7",X"25",X"13",X"27",X"06",X"7C",X"00",X"B2",X"7E",X"EB",X"91",X"BD",
		X"EC",X"28",X"6D",X"00",X"01",X"39",X"7A",X"00",X"B2",X"08",X"A6",X"00",X"DE",X"88",X"A6",X"00",
		X"08",X"DF",X"88",X"97",X"B8",X"CE",X"ED",X"5A",X"DF",X"AD",X"39",X"00",X"00",X"55",X"55",X"AA",
		X"55",X"5A",X"5A",X"96",X"69",X"66",X"66",X"CC",X"33",X"3C",X"3C",X"0F",X"F0",X"0D",X"20",X"0C",
		X"30",X"40",X"00",X"02",X"FF",X"00",X"FE",X"FE",X"80",X"30",X"63",X"05",X"2F",X"E0",X"67",X"F2",
		X"80",X"30",X"02",X"FE",X"00",X"FE",X"FE",X"00",X"02",X"FE",X"00",X"FE",X"FE",X"00",X"02",X"FE",
		X"00",X"FE",X"FE",X"00",X"06",X"FD",X"3F",X"00",X"FB",X"31",X"00",X"00",X"02",X"80",X"31",X"20",
		X"06",X"60",X"DE",X"70",X"D7",X"2A",X"21",X"00",X"01",X"2A",X"F0",X"01",X"1F",X"EB",X"01",X"19",
		X"F5",X"70",X"F3",X"0F",X"28",X"0E",X"28",X"0D",X"28",X"0C",X"28",X"0B",X"28",X"0A",X"28",X"09",
		X"28",X"08",X"28",X"40",X"10",X"0F",X"08",X"06",X"04",X"02",X"29",X"10",X"08",X"F8",X"22",X"10",
		X"0C",X"00",X"FA",X"23",X"10",X"0C",X"FC",X"00",X"23",X"10",X"07",X"FC",X"FC",X"FE",X"29",X"10",
		X"0E",X"00",X"FE",X"FA",X"26",X"3C",X"07",X"FC",X"70",X"DA",X"0F",X"08",X"0B",X"28",X"0D",X"00",
		X"FD",X"0C",X"28",X"0B",X"00",X"FD",X"0D",X"28",X"0C",X"00",X"FD",X"70",X"EF",X"10",X"01",X"02",
		X"2F",X"10",X"02",X"02",X"2F",X"10",X"04",X"02",X"2F",X"10",X"09",X"02",X"FE",X"2F",X"10",X"02",
		X"FE",X"2F",X"10",X"04",X"FE",X"2F",X"10",X"09",X"FE",X"00",X"2F",X"10",X"02",X"00",X"2F",X"10",
		X"04",X"00",X"2F",X"50",X"70",X"D7",X"0C",X"28",X"67",X"04",X"67",X"07",X"70",X"FA",X"63",X"00",
		X"38",X"37",X"40",X"63",X"00",X"36",X"39",X"40",X"10",X"FF",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"2F",X"2F",X"50",X"10",X"80",X"FE",X"2F",X"10",X"40",X"FE",X"2F",X"10",X"A0",X"00",
		X"FE",X"2F",X"10",X"50",X"00",X"FE",X"2F",X"10",X"28",X"00",X"FE",X"2F",X"10",X"14",X"00",X"FE",
		X"2F",X"10",X"0A",X"00",X"FE",X"2F",X"10",X"05",X"00",X"FE",X"2F",X"10",X"02",X"00",X"2F",X"10",
		X"01",X"00",X"2F",X"70",X"C3",X"53",X"80",X"10",X"8B",X"08",X"06",X"04",X"02",X"69",X"28",X"10",
		X"80",X"F8",X"62",X"23",X"10",X"88",X"00",X"FA",X"63",X"1D",X"10",X"88",X"FC",X"00",X"63",X"17",
		X"10",X"0B",X"FC",X"FC",X"FE",X"69",X"10",X"10",X"8A",X"00",X"FE",X"FA",X"66",X"09",X"3C",X"07",
		X"FC",X"70",X"D4",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"20",X"40",X"10",
		X"0F",X"02",X"FE",X"02",X"FE",X"2F",X"70",X"FD",X"10",X"74",X"02",X"02",X"02",X"02",X"2F",X"10",
		X"24",X"FE",X"FE",X"2F",X"10",X"50",X"FE",X"FE",X"2F",X"10",X"24",X"02",X"02",X"2F",X"70",X"E8",
		X"3C",X"81",X"70",X"FD",X"37",X"2F",X"00",X"01",X"37",X"F5",X"01",X"2D",X"F5",X"01",X"46",X"FA",
		X"70",X"F5",X"00",X"FA",X"20",X"80",X"F4",X"80",X"32",X"60",X"08",X"10",X"06",X"60",X"04",X"10",
		X"FA",X"70",X"F6",X"01",X"32",X"69",X"EB",X"01",X"28",X"6B",X"E7",X"01",X"20",X"6E",X"E3",X"80",
		X"19",X"69",X"00",X"10",X"04",X"01",X"19",X"20",X"64",X"88",X"01",X"20",X"20",X"96",X"B0",X"80",
		X"32",X"20",X"50",X"C7",X"20",X"AA",X"D1",X"21",X"FE",X"D0",X"80",X"ED",X"F3",X"EF",X"14",X"EE",
		X"04",X"EF",X"10",X"EE",X"2A",X"ED",X"E5",X"EE",X"3D",X"ED",X"E5",X"EE",X"66",X"EF",X"14",X"EE",
		X"78",X"EF",X"14",X"EE",X"B5",X"EF",X"10",X"EE",X"EF",X"EF",X"28",X"EE",X"F8",X"EF",X"40",X"EE",
		X"B5",X"EF",X"50",X"ED",X"AD",X"ED",X"DE",X"5F",X"D7",X"8D",X"48",X"48",X"8B",X"5B",X"C9",X"EF",
		X"D7",X"8A",X"97",X"8B",X"DE",X"8A",X"EE",X"00",X"DF",X"88",X"DE",X"8A",X"EE",X"02",X"E6",X"00",
		X"D7",X"8C",X"08",X"DF",X"8A",X"CE",X"ED",X"9B",X"DF",X"8E",X"7E",X"E9",X"D1",X"CC",X"38",X"3F",
		X"05",X"FC",X"00",X"29",X"07",X"1E",X"38",X"04",X"05",X"55",X"00",X"29",X"07",X"1E",X"38",X"0D",
		X"04",X"C0",X"00",X"29",X"07",X"1E",X"38",X"04",X"05",X"55",X"00",X"29",X"07",X"1E",X"38",X"3F",
		X"05",X"FC",X"00",X"29",X"07",X"1E",X"38",X"04",X"05",X"55",X"00",X"29",X"07",X"1E",X"38",X"0D",
		X"04",X"C0",X"00",X"29",X"07",X"1E",X"38",X"04",X"05",X"55",X"00",X"29",X"07",X"1E",X"38",X"3F",
		X"05",X"FC",X"00",X"29",X"07",X"1E",X"38",X"04",X"05",X"55",X"00",X"29",X"07",X"1E",X"38",X"0D",
		X"04",X"C0",X"00",X"29",X"07",X"1E",X"38",X"04",X"07",X"1C",X"00",X"29",X"07",X"1E",X"38",X"0D",
		X"04",X"C0",X"00",X"29",X"07",X"1E",X"38",X"29",X"07",X"1E",X"00",X"29",X"07",X"1E",X"38",X"37",
		X"03",X"2B",X"00",X"29",X"07",X"1E",X"38",X"3F",X"02",X"FE",X"00",X"29",X"07",X"1E",X"38",X"37",
		X"03",X"2B",X"00",X"29",X"07",X"1E",X"38",X"29",X"07",X"1E",X"00",X"29",X"07",X"1E",X"38",X"37",
		X"03",X"2B",X"00",X"29",X"07",X"1E",X"38",X"3F",X"02",X"FE",X"00",X"29",X"07",X"1E",X"38",X"37",
		X"03",X"2B",X"00",X"29",X"07",X"1E",X"38",X"29",X"07",X"1E",X"00",X"29",X"07",X"1E",X"38",X"37",
		X"03",X"2B",X"00",X"29",X"07",X"1E",X"38",X"3F",X"02",X"FE",X"00",X"29",X"07",X"1E",X"38",X"37",
		X"04",X"3A",X"00",X"29",X"07",X"1E",X"38",X"3F",X"02",X"FE",X"4F",X"7F",X"00",X"93",X"97",X"87",
		X"CE",X"EF",X"AD",X"A6",X"00",X"27",X"2D",X"7A",X"00",X"87",X"20",X"06",X"4C",X"BD",X"F1",X"1A",
		X"20",X"F1",X"08",X"DF",X"8E",X"BD",X"F1",X"1A",X"DF",X"8C",X"DE",X"8E",X"A6",X"00",X"97",X"96",
		X"A6",X"01",X"EE",X"02",X"DF",X"94",X"8D",X"0D",X"DE",X"8E",X"08",X"08",X"08",X"08",X"DF",X"8E",
		X"9C",X"8C",X"26",X"E8",X"39",X"CE",X"00",X"97",X"81",X"00",X"27",X"15",X"81",X"03",X"27",X"09",
		X"C6",X"01",X"E7",X"00",X"08",X"80",X"02",X"20",X"EF",X"C6",X"91",X"E7",X"00",X"6F",X"01",X"08",
		X"08",X"C6",X"7E",X"E7",X"00",X"C6",X"F0",X"E7",X"01",X"C6",X"DF",X"E7",X"02",X"DE",X"94",X"4F",
		X"F6",X"00",X"88",X"5C",X"D7",X"88",X"D4",X"96",X"54",X"89",X"00",X"54",X"89",X"00",X"54",X"89",
		X"00",X"54",X"89",X"00",X"54",X"89",X"00",X"54",X"89",X"00",X"54",X"89",X"00",X"48",X"48",X"48",
		X"48",X"48",X"B7",X"20",X"02",X"09",X"27",X"03",X"7E",X"00",X"97",X"39",X"96",X"81",X"44",X"98",
		X"81",X"44",X"44",X"76",X"00",X"80",X"76",X"00",X"81",X"39",X"DF",X"8C",X"9B",X"8D",X"97",X"8D",
		X"96",X"8C",X"89",X"00",X"97",X"8C",X"DE",X"8C",X"39",X"C6",X"BF",X"4F",X"B7",X"20",X"02",X"17",
		X"4A",X"26",X"FD",X"17",X"43",X"B7",X"20",X"02",X"8D",X"D2",X"4A",X"26",X"FD",X"5A",X"26",X"EB",
		X"39",X"C6",X"FF",X"7F",X"20",X"02",X"BD",X"F1",X"0C",X"96",X"81",X"20",X"00",X"4A",X"26",X"FB",
		X"73",X"20",X"02",X"C5",X"01",X"26",X"03",X"7A",X"20",X"02",X"17",X"4A",X"26",X"FD",X"73",X"20",
		X"02",X"5A",X"26",X"E2",X"39",X"C6",X"01",X"7F",X"20",X"02",X"BD",X"F1",X"0C",X"96",X"81",X"20",
		X"00",X"4A",X"26",X"FB",X"73",X"20",X"02",X"C5",X"01",X"26",X"03",X"7A",X"20",X"02",X"17",X"4A",
		X"26",X"FD",X"73",X"20",X"02",X"5C",X"26",X"E2",X"39",X"01",X"03",X"FF",X"80",X"FF",X"00",X"CE",
		X"F1",X"89",X"BD",X"E8",X"2A",X"7E",X"E8",X"43",X"48",X"03",X"01",X"0C",X"FF",X"00",X"86",X"FF",
		X"97",X"89",X"CE",X"F1",X"98",X"8D",X"EB",X"8D",X"02",X"20",X"FA",X"96",X"89",X"80",X"08",X"2A",
		X"03",X"97",X"89",X"39",X"32",X"32",X"39",X"C6",X"11",X"D7",X"AF",X"86",X"FE",X"97",X"94",X"86",
		X"9F",X"D6",X"AF",X"CE",X"01",X"C0",X"09",X"27",X"20",X"F7",X"00",X"93",X"B7",X"20",X"02",X"09",
		X"27",X"17",X"7A",X"00",X"93",X"26",X"F8",X"09",X"27",X"0F",X"D7",X"93",X"73",X"20",X"02",X"09",
		X"27",X"07",X"7A",X"00",X"93",X"26",X"F8",X"20",X"DD",X"D0",X"94",X"C1",X"10",X"22",X"D4",X"39",
		X"4F",X"B7",X"20",X"02",X"97",X"87",X"4F",X"91",X"87",X"26",X"03",X"73",X"20",X"02",X"C6",X"12",
		X"5A",X"26",X"FD",X"4C",X"2A",X"F1",X"73",X"20",X"02",X"7C",X"00",X"87",X"2A",X"E8",X"39",X"CE",
		X"00",X"93",X"6F",X"00",X"08",X"8C",X"00",X"A3",X"26",X"F8",X"86",X"18",X"97",X"93",X"CE",X"00",
		X"93",X"86",X"C0",X"97",X"87",X"5F",X"A6",X"01",X"AB",X"00",X"A7",X"01",X"2A",X"02",X"DB",X"87",
		X"74",X"00",X"87",X"08",X"08",X"8C",X"00",X"A3",X"26",X"EC",X"F7",X"20",X"02",X"7C",X"00",X"88",
		X"26",X"DC",X"CE",X"00",X"93",X"5F",X"A6",X"00",X"27",X"0B",X"81",X"37",X"26",X"04",X"C6",X"19",
		X"E7",X"02",X"6A",X"00",X"5C",X"08",X"08",X"8C",X"00",X"A3",X"26",X"EA",X"5D",X"26",X"BF",X"39",
		X"86",X"20",X"97",X"95",X"97",X"98",X"86",X"01",X"CE",X"00",X"01",X"C6",X"FF",X"97",X"93",X"DF",
		X"96",X"D7",X"94",X"D6",X"95",X"96",X"81",X"44",X"44",X"44",X"98",X"81",X"44",X"76",X"00",X"80",
		X"76",X"00",X"81",X"86",X"00",X"24",X"02",X"96",X"94",X"B7",X"20",X"02",X"DE",X"96",X"09",X"26",
		X"FD",X"5A",X"26",X"E1",X"D6",X"94",X"D0",X"93",X"27",X"09",X"DE",X"96",X"08",X"96",X"98",X"27",
		X"D0",X"20",X"CC",X"39",X"86",X"00",X"B7",X"20",X"02",X"CE",X"00",X"30",X"C6",X"25",X"5A",X"26",
		X"FD",X"73",X"20",X"02",X"09",X"26",X"F5",X"8B",X"10",X"2A",X"EB",X"20",X"E7",X"8D",X"09",X"7E",
		X"E1",X"46",X"86",X"17",X"8D",X"F7",X"20",X"FA",X"16",X"58",X"1B",X"1B",X"1B",X"CE",X"F3",X"2E",
		X"BD",X"F1",X"1A",X"A6",X"00",X"16",X"84",X"0F",X"97",X"95",X"54",X"54",X"54",X"54",X"D7",X"94",
		X"A6",X"01",X"16",X"54",X"54",X"54",X"54",X"D7",X"96",X"84",X"0F",X"97",X"87",X"DF",X"8A",X"CE",
		X"E2",X"25",X"7A",X"00",X"87",X"2B",X"08",X"A6",X"00",X"4C",X"BD",X"F1",X"1A",X"20",X"F3",X"DF",
		X"99",X"BD",X"E1",X"D0",X"DE",X"8A",X"A6",X"02",X"97",X"9B",X"BD",X"E1",X"E2",X"DE",X"8A",X"A6",
		X"03",X"97",X"97",X"A6",X"04",X"97",X"98",X"A6",X"05",X"16",X"A6",X"06",X"CE",X"F3",X"D6",X"BD",
		X"F1",X"1A",X"17",X"DF",X"9C",X"7F",X"00",X"A4",X"BD",X"F1",X"1A",X"DF",X"9E",X"39",X"81",X"24",
		X"00",X"00",X"00",X"16",X"31",X"41",X"45",X"00",X"00",X"00",X"0F",X"5B",X"F4",X"12",X"00",X"00",
		X"00",X"14",X"47",X"21",X"35",X"11",X"FF",X"00",X"0D",X"1B",X"F6",X"53",X"00",X"00",X"02",X"06",
		X"94",X"E3",X"12",X"00",X"00",X"02",X"06",X"9A",X"16",X"17",X"00",X"00",X"00",X"0A",X"10",X"41",
		X"02",X"D0",X"00",X"00",X"27",X"6D",X"FE",X"1A",X"00",X"00",X"00",X"08",X"6E",X"82",X"22",X"00",
		X"00",X"00",X"18",X"C6",X"51",X"3C",X"7F",X"00",X"00",X"0D",X"1B",X"B2",X"10",X"00",X"00",X"00",
		X"14",X"A4",X"FF",X"1F",X"14",X"01",X"01",X"04",X"1C",X"1C",X"1F",X"00",X"FF",X"FF",X"08",X"88",
		X"3D",X"5C",X"01",X"01",X"01",X"02",X"01",X"F4",X"15",X"00",X"00",X"00",X"08",X"1B",X"72",X"28",
		X"03",X"00",X"02",X"07",X"9A",X"D1",X"12",X"00",X"00",X"00",X"0C",X"00",X"3F",X"1F",X"11",X"01",
		X"07",X"04",X"1C",X"1F",X"F6",X"FE",X"FE",X"FE",X"01",X"21",X"01",X"17",X"00",X"00",X"00",X"08",
		X"1E",X"FF",X"16",X"00",X"00",X"00",X"08",X"88",X"F1",X"05",X"05",X"FF",X"01",X"20",X"0D",X"21",
		X"30",X"08",X"FF",X"01",X"27",X"0D",X"A0",X"98",X"90",X"88",X"80",X"78",X"70",X"68",X"60",X"58",
		X"50",X"44",X"40",X"01",X"01",X"02",X"02",X"04",X"04",X"08",X"08",X"10",X"10",X"30",X"60",X"C0",
		X"E0",X"01",X"01",X"02",X"02",X"03",X"04",X"05",X"06",X"07",X"08",X"09",X"0A",X"0C",X"80",X"7C",
		X"78",X"74",X"70",X"74",X"78",X"7C",X"80",X"01",X"01",X"02",X"02",X"04",X"04",X"08",X"08",X"10",
		X"20",X"28",X"30",X"38",X"40",X"48",X"50",X"60",X"70",X"80",X"A0",X"B0",X"C0",X"08",X"40",X"08",
		X"40",X"08",X"40",X"08",X"40",X"08",X"40",X"08",X"40",X"08",X"40",X"08",X"40",X"08",X"40",X"08",
		X"40",X"01",X"02",X"04",X"08",X"09",X"0A",X"0B",X"0C",X"0E",X"0F",X"10",X"12",X"14",X"16",X"40",
		X"10",X"08",X"01",X"01",X"01",X"01",X"01",X"02",X"02",X"03",X"03",X"04",X"04",X"05",X"06",X"08",
		X"0A",X"0C",X"10",X"14",X"18",X"20",X"30",X"40",X"50",X"40",X"30",X"20",X"10",X"0C",X"0A",X"08",
		X"07",X"06",X"05",X"04",X"03",X"02",X"02",X"01",X"01",X"01",X"07",X"08",X"09",X"0A",X"0C",X"08",
		X"17",X"18",X"19",X"1A",X"1B",X"1C",X"00",X"00",X"00",X"00",X"08",X"80",X"10",X"78",X"18",X"70",
		X"20",X"60",X"28",X"58",X"30",X"50",X"40",X"48",X"00",X"01",X"08",X"10",X"01",X"08",X"10",X"01",
		X"08",X"10",X"01",X"08",X"10",X"01",X"08",X"10",X"01",X"08",X"10",X"00",X"10",X"20",X"40",X"10",
		X"20",X"40",X"10",X"20",X"40",X"10",X"20",X"40",X"10",X"20",X"40",X"10",X"20",X"40",X"10",X"20",
		X"40",X"10",X"20",X"40",X"00",X"01",X"40",X"02",X"42",X"03",X"43",X"04",X"44",X"05",X"45",X"06",
		X"46",X"07",X"47",X"08",X"48",X"09",X"49",X"0A",X"4A",X"0B",X"4B",X"00",X"01",X"02",X"03",X"04",
		X"05",X"06",X"07",X"08",X"18",X"19",X"CE",X"F5",X"13",X"86",X"34",X"B7",X"20",X"03",X"09",X"09",
		X"86",X"80",X"B7",X"20",X"02",X"08",X"08",X"A6",X"01",X"27",X"27",X"C6",X"03",X"5A",X"26",X"FD",
		X"7A",X"00",X"87",X"E6",X"00",X"FB",X"20",X"02",X"F7",X"20",X"02",X"4A",X"27",X"E7",X"C6",X"07",
		X"5A",X"26",X"FD",X"01",X"01",X"E6",X"00",X"FB",X"20",X"02",X"F7",X"20",X"02",X"4A",X"26",X"EE",
		X"20",X"D3",X"39",X"FD",X"06",X"04",X"01",X"00",X"03",X"03",X"0B",X"FE",X"02",X"02",X"01",X"FB",
		X"03",X"03",X"01",X"FB",X"06",X"01",X"01",X"FE",X"02",X"05",X"0C",X"FA",X"0D",X"07",X"0E",X"F8",
		X"0D",X"09",X"0D",X"F6",X"0E",X"0C",X"0D",X"F4",X"0E",X"0C",X"0E",X"F4",X"0E",X"0C",X"0E",X"F1",
		X"0C",X"0C",X"0F",X"F3",X"0D",X"0A",X"10",X"F2",X"0C",X"0B",X"09",X"02",X"01",X"0A",X"08",X"EF",
		X"0B",X"0A",X"13",X"EF",X"0B",X"0B",X"0C",X"00",X"05",X"07",X"06",X"ED",X"0A",X"14",X"0A",X"D3",
		X"03",X"2D",X"02",X"BB",X"02",X"1B",X"07",X"E8",X"04",X"2B",X"01",X"E0",X"05",X"17",X"09",X"E7",
		X"07",X"18",X"08",X"EA",X"0A",X"17",X"09",X"E8",X"07",X"15",X"09",X"F2",X"02",X"01",X"01",X"E7",
		X"08",X"12",X"0A",X"F3",X"06",X"10",X"07",X"EC",X"0A",X"0A",X"12",X"F6",X"06",X"08",X"05",X"F4",
		X"0D",X"11",X"0B",X"F1",X"08",X"11",X"06",X"F1",X"0A",X"0C",X"0E",X"F1",X"08",X"12",X"06",X"EC",
		X"09",X"13",X"09",X"EF",X"07",X"0E",X"09",X"F0",X"0A",X"11",X"08",X"EF",X"08",X"16",X"08",X"F1",
		X"09",X"07",X"07",X"F7",X"08",X"0C",X"0C",X"F6",X"0A",X"02",X"02",X"FA",X"02",X"06",X"03",X"FA",
		X"04",X"01",X"02",X"FF",X"02",X"0A",X"06",X"F9",X"02",X"0D",X"03",X"FB",X"03",X"02",X"02",X"F9",
		X"06",X"02",X"04",X"FE",X"01",X"02",X"01",X"FD",X"01",X"01",X"01",X"F8",X"08",X"0B",X"0C",X"FE",
		X"03",X"02",X"02",X"F6",X"10",X"0D",X"0F",X"F1",X"0E",X"0B",X"13",X"ED",X"0B",X"0E",X"06",X"FD",
		X"05",X"14",X"08",X"E7",X"09",X"11",X"06",X"EE",X"04",X"16",X"09",X"E7",X"09",X"18",X"07",X"E3",
		X"05",X"1B",X"07",X"E8",X"09",X"1A",X"07",X"DF",X"05",X"1C",X"07",X"E8",X"09",X"1B",X"07",X"E3",
		X"06",X"1D",X"07",X"E8",X"09",X"1B",X"07",X"DD",X"05",X"19",X"08",X"E6",X"08",X"19",X"07",X"E1",
		X"05",X"1B",X"07",X"E5",X"08",X"1B",X"07",X"E4",X"06",X"1A",X"07",X"E7",X"08",X"1A",X"07",X"E9",
		X"07",X"14",X"07",X"ED",X"06",X"18",X"06",X"E7",X"08",X"16",X"0A",X"F0",X"0D",X"14",X"0B",X"EA",
		X"0A",X"15",X"0A",X"ED",X"0B",X"12",X"0C",X"EA",X"0A",X"15",X"0A",X"ED",X"0B",X"13",X"0B",X"EC",
		X"0B",X"17",X"0A",X"EA",X"0A",X"13",X"0B",X"ED",X"0B",X"13",X"0B",X"E9",X"09",X"15",X"0A",X"ED",
		X"0B",X"13",X"0B",X"EB",X"0A",X"14",X"0A",X"EE",X"0B",X"12",X"0B",X"EC",X"0A",X"15",X"0A",X"EB",
		X"0A",X"13",X"0B",X"EB",X"0A",X"14",X"0A",X"EF",X"0B",X"12",X"0B",X"EB",X"0A",X"17",X"09",X"EC",
		X"0A",X"10",X"0C",X"EE",X"0B",X"16",X"09",X"EC",X"0A",X"10",X"0C",X"ED",X"0A",X"14",X"0A",X"EC",
		X"0A",X"11",X"0B",X"F0",X"0B",X"12",X"0A",X"EC",X"09",X"11",X"0A",X"F3",X"0B",X"0B",X"0B",X"F3",
		X"0A",X"11",X"09",X"EF",X"09",X"0C",X"0A",X"F8",X"0D",X"0D",X"09",X"F1",X"09",X"10",X"09",X"F4",
		X"0B",X"0B",X"0B",X"F5",X"0B",X"0E",X"09",X"F4",X"0B",X"0E",X"0A",X"F1",X"0A",X"0F",X"0A",X"F3",
		X"0C",X"11",X"0A",X"EF",X"0A",X"10",X"0A",X"F2",X"0B",X"11",X"0A",X"EF",X"0B",X"13",X"0A",X"EF",
		X"0B",X"13",X"0A",X"ED",X"0A",X"11",X"0B",X"EC",X"0A",X"13",X"0B",X"EB",X"0A",X"13",X"0B",X"EB",
		X"0A",X"13",X"0B",X"EB",X"0A",X"13",X"0B",X"ED",X"0B",X"14",X"0B",X"EA",X"0A",X"13",X"0B",X"ED",
		X"0B",X"15",X"0A",X"ED",X"0B",X"13",X"0B",X"EE",X"0B",X"11",X"0B",X"F1",X"0B",X"0C",X"0C",X"F6",
		X"0B",X"04",X"0D",X"FF",X"05",X"03",X"06",X"F9",X"09",X"09",X"08",X"F8",X"07",X"07",X"06",X"FD",
		X"05",X"05",X"06",X"F1",X"08",X"14",X"09",X"F0",X"0C",X"0F",X"0D",X"F0",X"0C",X"0D",X"09",X"FF",
		X"06",X"05",X"06",X"F6",X"07",X"04",X"05",X"F6",X"07",X"11",X"0A",X"F2",X"0C",X"0B",X"0F",X"F3",
		X"0B",X"03",X"01",X"FD",X"07",X"0E",X"0B",X"F6",X"10",X"0B",X"0C",X"F9",X"12",X"09",X"0F",X"F5",
		X"0A",X"00",X"01",X"FA",X"03",X"05",X"08",X"02",X"01",X"07",X"09",X"FC",X"15",X"0A",X"0B",X"F1",
		X"09",X"07",X"09",X"FD",X"05",X"06",X"09",X"FC",X"06",X"01",X"03",X"FE",X"01",X"05",X"01",X"F4",
		X"08",X"0D",X"0C",X"F7",X"10",X"0A",X"0D",X"F8",X"0F",X"07",X"10",X"F6",X"0A",X"01",X"06",X"FC",
		X"02",X"0D",X"0B",X"EF",X"0A",X"06",X"07",X"00",X"02",X"0E",X"09",X"EB",X"09",X"0E",X"07",X"FC",
		X"04",X"0E",X"07",X"EB",X"09",X"17",X"06",X"F1",X"06",X"14",X"07",X"EB",X"08",X"12",X"06",X"EB",
		X"05",X"17",X"08",X"E8",X"08",X"12",X"06",X"EE",X"05",X"16",X"08",X"E8",X"08",X"19",X"06",X"EC",
		X"07",X"18",X"07",X"EA",X"08",X"19",X"06",X"EA",X"07",X"19",X"07",X"EC",X"08",X"13",X"06",X"EE",
		X"06",X"16",X"07",X"EC",X"08",X"13",X"07",X"EE",X"06",X"0E",X"07",X"EF",X"06",X"0E",X"07",X"F2",
		X"07",X"0D",X"07",X"F7",X"08",X"06",X"08",X"F9",X"07",X"08",X"07",X"FE",X"02",X"01",X"02",X"F9",
		X"0B",X"0C",X"0B",X"EE",X"09",X"0E",X"0B",X"F6",X"0D",X"0F",X"09",X"F1",X"0A",X"0F",X"0A",X"F3",
		X"0C",X"10",X"0B",X"EF",X"0B",X"11",X"0B",X"ED",X"0A",X"11",X"0B",X"EE",X"0A",X"0F",X"0C",X"ED",
		X"0A",X"13",X"0A",X"F0",X"0B",X"0F",X"0C",X"EF",X"0B",X"12",X"0A",X"F2",X"0C",X"0F",X"0B",X"EF",
		X"0A",X"0F",X"0B",X"F1",X"0B",X"10",X"0B",X"EF",X"0A",X"0B",X"0D",X"F3",X"0B",X"0F",X"0A",X"F2",
		X"09",X"01",X"01",X"FF",X"01",X"0A",X"0C",X"F3",X"0A",X"0B",X"0A",X"FB",X"0F",X"09",X"09",X"F7",
		X"0A",X"06",X"0C",X"F8",X"0A",X"08",X"0C",X"F7",X"0B",X"0B",X"0A",X"F5",X"0B",X"0B",X"0B",X"F2",
		X"0A",X"10",X"0A",X"F2",X"0B",X"0D",X"0C",X"ED",X"09",X"10",X"0B",X"F0",X"0B",X"10",X"0B",X"EE",
		X"0A",X"11",X"0B",X"ED",X"0A",X"11",X"0B",X"EE",X"0A",X"0F",X"0C",X"EE",X"0A",X"10",X"0B",X"EE",
		X"0A",X"11",X"0B",X"ED",X"0A",X"11",X"0B",X"ED",X"0A",X"10",X"0C",X"ED",X"0A",X"13",X"0A",X"EF",
		X"0B",X"11",X"0B",X"EF",X"0B",X"11",X"0B",X"ED",X"0A",X"12",X"0B",X"EC",X"0A",X"12",X"0B",X"EF",
		X"0B",X"12",X"0A",X"EF",X"0B",X"11",X"0B",X"ED",X"0A",X"11",X"0B",X"EF",X"0B",X"11",X"0B",X"EE",
		X"0A",X"11",X"0B",X"ED",X"0A",X"11",X"0B",X"EF",X"0B",X"11",X"0B",X"ED",X"0A",X"11",X"0B",X"F0",
		X"0B",X"10",X"0B",X"EE",X"0A",X"10",X"0B",X"F0",X"0B",X"10",X"0B",X"EF",X"0A",X"0E",X"0C",X"F1",
		X"0B",X"0E",X"0B",X"F3",X"0B",X"0C",X"0B",X"F4",X"0B",X"0C",X"0B",X"F4",X"0B",X"0C",X"0B",X"F5",
		X"0B",X"0B",X"0B",X"F8",X"0D",X"09",X"0A",X"FA",X"0C",X"05",X"0B",X"FC",X"0B",X"00",X"03",X"FF",
		X"02",X"03",X"0A",X"FE",X"0A",X"00",X"02",X"FD",X"04",X"03",X"0A",X"FE",X"07",X"00",X"02",X"FF",
		X"07",X"04",X"09",X"FA",X"07",X"02",X"10",X"FA",X"09",X"09",X"09",X"F9",X"0A",X"05",X"10",X"F6",
		X"0B",X"09",X"0C",X"F7",X"09",X"08",X"08",X"F6",X"07",X"04",X"08",X"FF",X"05",X"08",X"09",X"EF",
		X"09",X"11",X"0A",X"F2",X"09",X"0C",X"08",X"F0",X"07",X"0B",X"09",X"F8",X"08",X"0D",X"07",X"EF",
		X"09",X"13",X"09",X"ED",X"08",X"13",X"08",X"EE",X"09",X"0E",X"09",X"F5",X"06",X"0A",X"08",X"EF",
		X"09",X"13",X"09",X"EC",X"08",X"12",X"09",X"ED",X"09",X"11",X"09",X"F0",X"06",X"0C",X"08",X"EF",
		X"09",X"13",X"09",X"EB",X"08",X"14",X"09",X"EB",X"09",X"12",X"09",X"EF",X"07",X"11",X"07",X"F0",
		X"09",X"11",X"09",X"F0",X"09",X"15",X"07",X"EE",X"09",X"12",X"09",X"F0",X"08",X"0D",X"08",X"EE",
		X"07",X"0F",X"09",X"F4",X"09",X"09",X"08",X"F6",X"08",X"0F",X"08",X"F1",X"09",X"0E",X"09",X"F3",
		X"08",X"09",X"08",X"F8",X"08",X"0B",X"08",X"F2",X"08",X"0E",X"09",X"F4",X"0A",X"0E",X"08",X"F4",
		X"08",X"08",X"08",X"FA",X"09",X"08",X"08",X"F6",X"08",X"0B",X"09",X"F2",X"08",X"0C",X"09",X"F5",
		X"09",X"0C",X"08",X"F6",X"08",X"0A",X"08",X"F1",X"07",X"0E",X"09",X"F1",X"09",X"0F",X"09",X"F0",
		X"08",X"0B",X"09",X"F5",X"07",X"0B",X"08",X"F2",X"08",X"0C",X"09",X"F7",X"09",X"07",X"09",X"F8",
		X"08",X"08",X"09",X"F9",X"09",X"05",X"0A",X"FB",X"07",X"02",X"02",X"FE",X"01",X"03",X"06",X"FD",
		X"07",X"07",X"08",X"F6",X"09",X"08",X"0A",X"FA",X"0A",X"04",X"0A",X"FE",X"07",X"00",X"01",X"FF",
		X"04",X"02",X"0A",X"FC",X"0A",X"06",X"09",X"FA",X"08",X"03",X"08",X"FE",X"07",X"03",X"07",X"FD",
		X"0B",X"07",X"08",X"F7",X"09",X"09",X"09",X"F8",X"08",X"06",X"09",X"FB",X"0B",X"08",X"08",X"F9",
		X"09",X"06",X"08",X"FA",X"07",X"06",X"08",X"FB",X"0A",X"05",X"0B",X"F9",X"09",X"07",X"09",X"F8",
		X"08",X"06",X"0A",X"FC",X"0B",X"04",X"0A",X"FE",X"0A",X"FE",X"03",X"FF",X"08",X"05",X"08",X"F9",
		X"0A",X"07",X"09",X"FC",X"09",X"04",X"08",X"FD",X"0C",X"03",X"08",X"FF",X"06",X"02",X"07",X"FA",
		X"08",X"08",X"09",X"F6",X"08",X"08",X"0A",X"FA",X"09",X"01",X"09",X"05",X"01",X"00",X"03",X"01",
		X"01",X"03",X"08",X"FB",X"0B",X"08",X"08",X"F8",X"08",X"06",X"0A",X"FB",X"09",X"02",X"06",X"FE",
		X"05",X"05",X"0B",X"F8",X"0A",X"07",X"09",X"FA",X"07",X"06",X"09",X"F9",X"0A",X"06",X"08",X"FB",
		X"07",X"06",X"09",X"F8",X"08",X"04",X"09",X"FD",X"07",X"04",X"0A",X"FD",X"08",X"02",X"02",X"FC",
		X"03",X"01",X"01",X"FB",X"04",X"05",X"0B",X"FC",X"09",X"05",X"07",X"F8",X"08",X"07",X"0A",X"FB",
		X"09",X"06",X"08",X"F9",X"0A",X"06",X"09",X"FD",X"08",X"01",X"07",X"00",X"02",X"02",X"03",X"FF",
		X"02",X"02",X"03",X"FE",X"0C",X"03",X"0D",X"FB",X"0B",X"06",X"0A",X"FA",X"0C",X"08",X"0A",X"F8",
		X"0A",X"07",X"09",X"FB",X"06",X"05",X"07",X"F9",X"0B",X"0B",X"09",X"F7",X"09",X"05",X"0A",X"FA",
		X"09",X"0B",X"09",X"F3",X"0A",X"0A",X"0B",X"FB",X"0D",X"02",X"18",X"F8",X"09",X"07",X"0C",X"FB",
		X"08",X"00",X"02",X"FF",X"02",X"02",X"02",X"FC",X"07",X"04",X"10",X"F7",X"09",X"06",X"0A",X"FF",
		X"06",X"00",X"02",X"FF",X"02",X"00",X"02",X"FC",X"09",X"03",X"10",X"FC",X"0C",X"04",X"0D",X"FD",
		X"0B",X"00",X"03",X"FE",X"02",X"04",X"01",X"FF",X"04",X"03",X"0C",X"FB",X"08",X"02",X"08",X"FF",
		X"03",X"00",X"01",X"FF",X"03",X"04",X"08",X"FB",X"0A",X"03",X"0E",X"00",X"02",X"00",X"01",X"FD",
		X"0A",X"02",X"0B",X"00",X"02",X"01",X"02",X"FF",X"02",X"01",X"03",X"FE",X"0E",X"04",X"0C",X"FA",
		X"0A",X"05",X"09",X"FD",X"08",X"03",X"06",X"FE",X"0A",X"01",X"03",X"00",X"01",X"01",X"0C",X"FE",
		X"09",X"03",X"08",X"FE",X"09",X"01",X"07",X"FF",X"09",X"01",X"0B",X"FF",X"0B",X"03",X"09",X"FC",
		X"09",X"04",X"09",X"FD",X"0A",X"03",X"09",X"FE",X"0C",X"01",X"0A",X"00",X"06",X"FD",X"01",X"FF",
		X"02",X"02",X"08",X"FE",X"0B",X"02",X"0A",X"FE",X"08",X"01",X"07",X"00",X"02",X"01",X"01",X"FF",
		X"08",X"01",X"02",X"FF",X"02",X"01",X"03",X"00",X"03",X"00",X"02",X"FC",X"01",X"01",X"03",X"00",
		X"02",X"01",X"0B",X"FE",X"0B",X"03",X"08",X"FF",X"08",X"FE",X"01",X"00",X"06",X"FF",X"02",X"00",
		X"06",X"00",X"0B",X"00",X"07",X"02",X"03",X"00",X"0B",X"00",X"00",X"7F",X"20",X"00",X"86",X"FF",
		X"97",X"94",X"CE",X"FB",X"8E",X"DF",X"95",X"DE",X"95",X"A6",X"00",X"27",X"2B",X"97",X"93",X"E6",
		X"01",X"08",X"08",X"DF",X"95",X"96",X"94",X"B7",X"20",X"02",X"96",X"93",X"CE",X"00",X"06",X"09",
		X"26",X"FD",X"4A",X"26",X"F7",X"7F",X"20",X"02",X"96",X"93",X"CE",X"00",X"06",X"09",X"26",X"FD",
		X"4A",X"26",X"F7",X"5A",X"26",X"DF",X"20",X"CF",X"86",X"80",X"B7",X"20",X"00",X"39",X"01",X"30",
		X"02",X"0C",X"03",X"08",X"04",X"08",X"06",X"08",X"08",X"04",X"0C",X"04",X"10",X"04",X"20",X"02",
		X"40",X"01",X"60",X"01",X"80",X"01",X"A0",X"01",X"C0",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"2E",X"E0",X"01",X"E0",X"43",X"E0",X"01");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
