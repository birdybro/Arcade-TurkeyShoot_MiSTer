library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity turkey_shoot_graph1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of turkey_shoot_graph1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"FF",X"FF",X"EF",
		X"22",X"FF",X"F2",X"22",X"22",X"FA",X"22",X"C2",X"EE",X"2A",X"EE",X"EE",X"DD",X"AA",X"2E",X"DE",
		X"CC",X"AF",X"2A",X"CE",X"EE",X"CC",X"AE",X"EE",X"AA",X"CC",X"AA",X"AA",X"77",X"CC",X"F7",X"77",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"88",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"66",X"66",X"66",X"66",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"33",X"FF",X"FF",X"FF",X"F3",X"F3",X"3F",X"FF",X"F3",X"F3",X"F3",X"FF",X"F3",X"F3",X"F3",
		X"FF",X"F3",X"F3",X"F3",X"FF",X"3F",X"F3",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"11",
		X"FF",X"FF",X"FF",X"AF",X"FF",X"FF",X"FF",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"11",
		X"77",X"77",X"9F",X"77",X"77",X"77",X"9F",X"77",X"77",X"77",X"9F",X"77",X"77",X"77",X"9F",X"77",
		X"77",X"77",X"9F",X"77",X"77",X"77",X"9F",X"77",X"77",X"77",X"9F",X"77",X"77",X"77",X"9F",X"77",
		X"77",X"77",X"9F",X"77",X"77",X"77",X"9F",X"77",X"77",X"77",X"9F",X"77",X"77",X"77",X"9F",X"77",
		X"77",X"77",X"9F",X"77",X"77",X"77",X"9F",X"77",X"FF",X"FF",X"9F",X"FF",X"77",X"77",X"9F",X"77",
		X"77",X"FF",X"77",X"FF",X"99",X"FF",X"99",X"FC",X"88",X"CF",X"88",X"C8",X"27",X"57",X"57",X"57",
		X"27",X"57",X"C7",X"57",X"27",X"57",X"57",X"57",X"27",X"C5",X"C7",X"57",X"88",X"88",X"88",X"88",
		X"99",X"99",X"99",X"99",X"88",X"88",X"88",X"88",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",X"C7",
		X"27",X"27",X"27",X"27",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",
		X"F7",X"77",X"77",X"FF",X"99",X"99",X"F9",X"FF",X"88",X"8F",X"88",X"88",X"55",X"25",X"5F",X"25",
		X"52",X"25",X"25",X"25",X"55",X"25",X"55",X"25",X"55",X"25",X"25",X"25",X"88",X"88",X"88",X"F8",
		X"99",X"99",X"99",X"FC",X"88",X"88",X"88",X"C8",X"CC",X"CC",X"CF",X"6C",X"CC",X"CC",X"CF",X"CF",
		X"22",X"22",X"2F",X"2F",X"22",X"22",X"2F",X"2F",X"22",X"22",X"2F",X"2F",X"22",X"22",X"2F",X"2F",
		X"DF",X"FF",X"FF",X"FF",X"DD",X"FF",X"FF",X"DD",X"FF",X"DD",X"DD",X"FF",X"FF",X"FF",X"FF",X"DD",
		X"EE",X"FF",X"DF",X"3D",X"FE",X"DD",X"33",X"F3",X"DD",X"D3",X"FF",X"FF",X"FD",X"E3",X"F1",X"1F",
		X"FF",X"D3",X"F1",X"1F",X"FD",X"E3",X"F1",X"1F",X"EE",X"D3",X"11",X"1F",X"EE",X"D3",X"F1",X"1F",
		X"EE",X"D3",X"F1",X"1F",X"DD",X"D3",X"F1",X"FF",X"FF",X"D3",X"FF",X"3F",X"FF",X"EE",X"33",X"F3",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"DD",X"DD",X"FF",X"FF",
		X"D3",X"FD",X"33",X"FF",X"3F",X"33",X"FF",X"FF",X"F1",X"FF",X"11",X"FF",X"F1",X"F1",X"FF",X"FF",
		X"F1",X"1F",X"FF",X"FF",X"F1",X"1F",X"11",X"DF",X"F1",X"1F",X"FF",X"DD",X"F1",X"1F",X"FF",X"ED",
		X"F1",X"1F",X"11",X"DD",X"FF",X"F1",X"FF",X"DD",X"F3",X"FF",X"33",X"DD",X"3D",X"33",X"DD",X"DD",
		X"F7",X"77",X"77",X"7B",X"F7",X"B1",X"B1",X"B1",X"F1",X"22",X"22",X"22",X"B2",X"21",X"22",X"11",
		X"12",X"F2",X"F1",X"1F",X"B2",X"22",X"21",X"11",X"12",X"12",X"21",X"1F",X"B2",X"2F",X"21",X"1F",
		X"12",X"F2",X"22",X"2F",X"B2",X"22",X"22",X"22",X"F1",X"22",X"22",X"22",X"F7",X"B1",X"B1",X"B1",
		X"F7",X"FF",X"FF",X"FF",X"F9",X"FF",X"AA",X"AA",X"F9",X"7F",X"CC",X"CC",X"F9",X"77",X"CC",X"CC",
		X"22",X"77",X"77",X"78",X"22",X"B1",X"B1",X"B1",X"22",X"22",X"22",X"22",X"21",X"12",X"21",X"11",
		X"21",X"1F",X"21",X"FF",X"21",X"1F",X"F1",X"11",X"21",X"1F",X"F1",X"F1",X"21",X"1F",X"F1",X"F2",
		X"22",X"2F",X"22",X"F2",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"B1",X"B1",X"B1",X"B1",
		X"77",X"FF",X"FF",X"77",X"77",X"AA",X"AA",X"77",X"99",X"AC",X"AC",X"99",X"99",X"AC",X"AC",X"99",
		X"76",X"72",X"CC",X"22",X"7F",X"72",X"00",X"C2",X"77",X"72",X"CA",X"02",X"77",X"72",X"2A",X"C2",
		X"77",X"72",X"00",X"22",X"77",X"72",X"0A",X"CC",X"77",X"72",X"C0",X"00",X"76",X"00",X"CA",X"CC",
		X"76",X"87",X"44",X"77",X"7F",X"72",X"CA",X"44",X"77",X"72",X"2A",X"CC",X"77",X"72",X"44",X"2C",
		X"77",X"72",X"4A",X"2C",X"77",X"7C",X"C4",X"CC",X"77",X"44",X"2A",X"44",X"76",X"72",X"2A",X"CC",
		X"F1",X"11",X"F7",X"77",X"F1",X"1F",X"F7",X"70",X"F1",X"1F",X"77",X"70",X"F1",X"1F",X"07",X"70",
		X"F1",X"1F",X"07",X"70",X"F1",X"11",X"07",X"70",X"FF",X"FF",X"07",X"70",X"4F",X"F4",X"07",X"70",
		X"F4",X"F4",X"07",X"70",X"F4",X"F4",X"07",X"70",X"F4",X"74",X"07",X"70",X"47",X"74",X"07",X"70",
		X"88",X"70",X"07",X"70",X"78",X"70",X"07",X"70",X"88",X"A0",X"07",X"70",X"22",X"7F",X"F2",X"2F",
		X"FF",X"00",X"FF",X"FF",X"FF",X"F4",X"FF",X"FF",X"F0",X"11",X"FF",X"FF",X"F0",X"F4",X"FF",X"FF",
		X"F0",X"F4",X"FF",X"FF",X"F0",X"11",X"FF",X"FF",X"F0",X"F4",X"FF",X"FF",X"F0",X"F4",X"FF",X"FF",
		X"F0",X"F4",X"FF",X"FF",X"F0",X"11",X"FF",X"FF",X"FF",X"F4",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"FF",X"FF",X"FF",X"99",X"FF",X"FF",X"FF",X"99",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",
		X"79",X"AA",X"AA",X"AA",X"79",X"AC",X"CA",X"CC",X"79",X"AC",X"2A",X"2C",X"79",X"A2",X"2A",X"32",
		X"79",X"A2",X"2A",X"32",X"79",X"A2",X"2A",X"32",X"79",X"A2",X"2A",X"32",X"79",X"A2",X"2A",X"32",
		X"79",X"A2",X"CA",X"3C",X"79",X"AC",X"CA",X"CC",X"88",X"88",X"00",X"08",X"8E",X"EE",X"EE",X"0E",
		X"8E",X"EE",X"00",X"0E",X"8E",X"EE",X"EE",X"E0",X"88",X"88",X"88",X"88",X"77",X"AA",X"AA",X"77",
		X"AA",X"AA",X"AA",X"AA",X"CC",X"CC",X"CC",X"CA",X"CC",X"C3",X"2C",X"2A",X"23",X"22",X"22",X"2A",
		X"32",X"22",X"C2",X"CA",X"22",X"22",X"C2",X"2A",X"2C",X"22",X"CC",X"CA",X"3C",X"22",X"C2",X"CA",
		X"C3",X"32",X"C2",X"CA",X"CC",X"CC",X"C2",X"CA",X"88",X"00",X"00",X"88",X"E0",X"0E",X"00",X"EE",
		X"E0",X"0E",X"EE",X"EE",X"E0",X"00",X"00",X"EE",X"88",X"88",X"88",X"88",X"AA",X"7A",X"AA",X"AA",
		X"FF",X"F9",X"FF",X"9F",X"FF",X"79",X"FF",X"91",X"FF",X"79",X"77",X"91",X"FF",X"17",X"71",X"91",
		X"FF",X"11",X"71",X"91",X"FF",X"11",X"71",X"97",X"FF",X"77",X"71",X"77",X"FF",X"11",X"99",X"99",
		X"FF",X"11",X"73",X"77",X"FF",X"19",X"93",X"99",X"FF",X"77",X"73",X"77",X"FF",X"99",X"99",X"99",
		X"FF",X"33",X"77",X"33",X"FF",X"99",X"99",X"39",X"FF",X"77",X"77",X"37",X"FF",X"33",X"33",X"37",
		X"CC",X"AC",X"CA",X"AA",X"CC",X"AC",X"CA",X"CC",X"44",X"A4",X"4A",X"44",X"44",X"A4",X"4A",X"44",
		X"44",X"A4",X"4A",X"44",X"44",X"A4",X"4A",X"44",X"44",X"A4",X"4A",X"44",X"44",X"A4",X"4A",X"AA",
		X"CC",X"AC",X"CA",X"44",X"CC",X"AC",X"CA",X"44",X"99",X"99",X"99",X"44",X"77",X"77",X"77",X"4C",
		X"77",X"77",X"77",X"CC",X"77",X"77",X"77",X"DD",X"88",X"88",X"88",X"CC",X"66",X"66",X"66",X"66",
		X"88",X"88",X"88",X"88",X"33",X"F3",X"77",X"B7",X"E3",X"23",X"22",X"BB",X"33",X"33",X"2B",X"BB",
		X"33",X"33",X"2B",X"BB",X"F3",X"33",X"2B",X"FB",X"F3",X"33",X"2B",X"AB",X"FF",X"3F",X"2F",X"A7",
		X"4F",X"3F",X"2A",X"F7",X"4F",X"F2",X"FC",X"BF",X"4F",X"F2",X"CC",X"BC",X"7F",X"F2",X"BF",X"BC",
		X"7F",X"F2",X"BB",X"BF",X"7F",X"FC",X"BB",X"F7",X"7F",X"CC",X"BB",X"77",X"7F",X"CF",X"FF",X"77",
		X"88",X"88",X"88",X"88",X"55",X"55",X"E7",X"77",X"55",X"55",X"74",X"4C",X"55",X"55",X"44",X"44",
		X"7F",X"5F",X"44",X"44",X"77",X"5F",X"4F",X"44",X"77",X"5C",X"7C",X"F4",X"77",X"5C",X"46",X"AF",
		X"77",X"5F",X"44",X"A7",X"77",X"5F",X"44",X"A7",X"77",X"5F",X"44",X"A7",X"77",X"5F",X"74",X"A7",
		X"77",X"5F",X"77",X"FF",X"77",X"5C",X"77",X"44",X"77",X"5C",X"77",X"D4",X"77",X"5F",X"77",X"44",
		X"AE",X"CF",X"CF",X"EE",X"77",X"CF",X"CF",X"77",X"77",X"CF",X"CF",X"77",X"77",X"CF",X"CF",X"88",
		X"78",X"CF",X"CF",X"88",X"78",X"CF",X"CF",X"88",X"78",X"CF",X"2F",X"88",X"78",X"CF",X"2F",X"88",
		X"78",X"2F",X"2F",X"88",X"FA",X"2F",X"2F",X"AE",X"78",X"2F",X"2F",X"88",X"78",X"2F",X"2F",X"88",
		X"78",X"2F",X"2F",X"88",X"78",X"2F",X"2F",X"88",X"AE",X"2F",X"2F",X"EE",X"76",X"2F",X"2F",X"66",
		X"CC",X"CA",X"AA",X"CA",X"CC",X"CA",X"CA",X"CA",X"22",X"2A",X"2A",X"2A",X"22",X"2A",X"2A",X"2A",
		X"22",X"2A",X"2A",X"2A",X"22",X"2A",X"2A",X"2A",X"22",X"2A",X"2A",X"2A",X"2C",X"2A",X"AA",X"2A",
		X"CC",X"CA",X"2A",X"CA",X"CC",X"CA",X"2A",X"CA",X"99",X"9A",X"2A",X"99",X"77",X"7A",X"CA",X"77",
		X"77",X"7A",X"CA",X"77",X"77",X"7A",X"AA",X"77",X"88",X"8C",X"CC",X"88",X"66",X"66",X"66",X"66",
		X"78",X"2F",X"2F",X"88",X"78",X"2F",X"2F",X"88",X"78",X"2F",X"2F",X"88",X"78",X"2F",X"2F",X"88",
		X"78",X"2F",X"2F",X"88",X"78",X"2F",X"2F",X"88",X"78",X"2F",X"2F",X"88",X"78",X"F2",X"F2",X"88",
		X"78",X"FF",X"FF",X"88",X"FA",X"2F",X"2F",X"AE",X"78",X"AA",X"DF",X"88",X"78",X"77",X"6F",X"88",
		X"78",X"77",X"6F",X"88",X"78",X"77",X"6F",X"88",X"78",X"CC",X"67",X"88",X"66",X"66",X"66",X"66",
		X"19",X"1E",X"77",X"E1",X"F1",X"7E",X"77",X"E1",X"F7",X"7E",X"11",X"11",X"F7",X"7E",X"77",X"E7",
		X"F7",X"44",X"77",X"E7",X"F7",X"4E",X"77",X"E7",X"F7",X"49",X"49",X"49",X"F7",X"47",X"74",X"74",
		X"44",X"4E",X"47",X"44",X"47",X"4E",X"77",X"E4",X"47",X"4E",X"77",X"E4",X"F4",X"7E",X"77",X"E4",
		X"F9",X"7E",X"44",X"44",X"FF",X"7E",X"77",X"E7",X"77",X"7E",X"77",X"E7",X"77",X"7E",X"77",X"E7",
		X"9F",X"22",X"22",X"F7",X"FF",X"22",X"22",X"F7",X"77",X"11",X"22",X"F7",X"77",X"22",X"2C",X"F7",
		X"79",X"2C",X"CC",X"F9",X"7F",X"EE",X"EE",X"FF",X"7F",X"44",X"77",X"99",X"44",X"77",X"77",X"77",
		X"7F",X"22",X"22",X"FF",X"77",X"44",X"22",X"F7",X"77",X"22",X"22",X"F7",X"77",X"22",X"22",X"F7",
		X"99",X"44",X"22",X"F7",X"FF",X"E2",X"22",X"F7",X"7F",X"22",X"22",X"F7",X"7F",X"22",X"22",X"F7",
		X"9F",X"22",X"22",X"F7",X"FF",X"22",X"22",X"F7",X"77",X"00",X"22",X"F7",X"00",X"22",X"2C",X"F7",
		X"79",X"2C",X"CC",X"F9",X"7F",X"00",X"EE",X"FF",X"7F",X"97",X"77",X"99",X"7F",X"77",X"77",X"77",
		X"7F",X"00",X"22",X"FF",X"77",X"22",X"22",X"F7",X"77",X"22",X"22",X"F7",X"77",X"22",X"22",X"F7",
		X"99",X"11",X"22",X"F7",X"11",X"E2",X"22",X"F7",X"7F",X"A2",X"22",X"F7",X"7F",X"11",X"22",X"F7",
		X"99",X"00",X"77",X"E7",X"FF",X"0E",X"77",X"E7",X"F7",X"0E",X"07",X"07",X"F7",X"0E",X"70",X"E0",
		X"00",X"0E",X"07",X"00",X"07",X"0E",X"77",X"E0",X"07",X"09",X"99",X"90",X"F0",X"77",X"77",X"70",
		X"F7",X"7E",X"00",X"07",X"F7",X"7E",X"77",X"E7",X"F7",X"11",X"77",X"E7",X"F7",X"1E",X"77",X"E7",
		X"F9",X"1E",X"17",X"17",X"FF",X"1E",X"71",X"A1",X"11",X"1E",X"17",X"11",X"17",X"1E",X"77",X"A1",
		X"77",X"8F",X"8F",X"FF",X"77",X"8F",X"7F",X"FF",X"AE",X"8F",X"66",X"66",X"FF",X"8F",X"37",X"77",
		X"EF",X"8F",X"73",X"37",X"CF",X"83",X"37",X"37",X"FC",X"83",X"37",X"37",X"FC",X"83",X"73",X"77",
		X"F7",X"83",X"77",X"77",X"F7",X"9F",X"33",X"33",X"F7",X"9F",X"8F",X"FF",X"F7",X"9F",X"8F",X"FF",
		X"F7",X"9F",X"DE",X"FF",X"FF",X"9D",X"DD",X"FF",X"FC",X"DD",X"DD",X"FF",X"F7",X"DD",X"DD",X"FF",
		X"44",X"44",X"33",X"F7",X"44",X"44",X"77",X"F7",X"44",X"44",X"77",X"F7",X"44",X"44",X"77",X"F7",
		X"44",X"44",X"33",X"F7",X"74",X"47",X"73",X"F7",X"74",X"47",X"33",X"F7",X"77",X"77",X"77",X"F7",
		X"77",X"44",X"33",X"F7",X"77",X"44",X"77",X"F7",X"77",X"47",X"77",X"F7",X"44",X"47",X"77",X"F7",
		X"44",X"47",X"33",X"F7",X"74",X"47",X"77",X"F7",X"FF",X"FF",X"07",X"FF",X"77",X"77",X"70",X"F7",
		X"88",X"FF",X"FF",X"FF",X"99",X"CC",X"FF",X"1F",X"99",X"77",X"FF",X"F1",X"99",X"77",X"FF",X"F1",
		X"99",X"79",X"99",X"71",X"99",X"78",X"88",X"71",X"99",X"F8",X"88",X"17",X"99",X"F8",X"FF",X"99",
		X"99",X"98",X"88",X"8F",X"99",X"88",X"88",X"1F",X"99",X"88",X"88",X"81",X"FF",X"FF",X"FF",X"FF",
		X"B8",X"8B",X"B8",X"88",X"B9",X"9B",X"B9",X"99",X"B8",X"8B",X"B8",X"88",X"FF",X"FF",X"FF",X"FF",
		X"11",X"11",X"11",X"11",X"C1",X"1C",X"C1",X"11",X"1C",X"11",X"1C",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"CC",X"CC",X"CC",X"CC",X"99",X"9F",X"99",X"99",X"88",X"8C",X"8F",X"8F",
		X"8F",X"88",X"8C",X"8F",X"F8",X"88",X"88",X"8F",X"C8",X"8F",X"88",X"8F",X"FF",X"FF",X"FF",X"FF",
		X"66",X"66",X"66",X"66",X"EE",X"67",X"66",X"66",X"6E",X"66",X"66",X"EE",X"66",X"66",X"66",X"66",
		X"FF",X"FF",X"FF",X"FF",X"77",X"77",X"77",X"77",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"11",X"11",X"11",X"CC",X"11",X"11",X"11",X"CC",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"C1",X"11",X"11",X"11",X"1C",X"11",
		X"C1",X"11",X"11",X"11",X"1C",X"11",X"C1",X"11",X"11",X"C1",X"1C",X"11",X"11",X"1C",X"11",X"11",
		X"BB",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"FF",X"1F",X"FB",X"FF",X"FF",X"FF",X"FF",X"BB",X"FF",
		X"FF",X"99",X"99",X"FF",X"FF",X"81",X"11",X"FF",X"99",X"81",X"18",X"77",X"88",X"81",X"18",X"17",
		X"88",X"81",X"11",X"17",X"88",X"81",X"11",X"17",X"18",X"88",X"18",X"77",X"FF",X"FF",X"FF",X"FF",
		X"B8",X"B8",X"88",X"8B",X"B9",X"B9",X"99",X"9B",X"B8",X"B8",X"88",X"8B",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"3F",X"3F",X"33",X"3F",X"FF",X"3F",X"3F",X"F3",X"FF",X"3F",X"33",X"F3",
		X"3F",X"3F",X"3F",X"F3",X"FF",X"3F",X"33",X"3F",X"FF",X"FF",X"FF",X"FF",X"1F",X"FF",X"FF",X"FF",
		X"F1",X"1F",X"FF",X"FF",X"11",X"1F",X"FF",X"FF",X"F1",X"FF",X"FF",X"FF",X"F1",X"1F",X"FF",X"FF",
		X"CC",X"FF",X"AA",X"FA",X"CC",X"F6",X"FA",X"FA",X"2C",X"F6",X"6C",X"F6",X"22",X"C7",X"FC",X"CF",
		X"22",X"F7",X"6C",X"FC",X"22",X"C7",X"FF",X"CF",X"22",X"F7",X"F6",X"FC",X"22",X"C7",X"FF",X"CF",
		X"22",X"F7",X"AF",X"EC",X"77",X"C7",X"FF",X"CF",X"77",X"FC",X"FE",X"FA",X"77",X"CF",X"CC",X"AA",
		X"77",X"FF",X"C2",X"AA",X"76",X"FF",X"AA",X"AA",X"66",X"FF",X"EA",X"2E",X"FF",X"FF",X"66",X"66",
		X"89",X"AA",X"CC",X"F8",X"89",X"EA",X"C2",X"F8",X"F8",X"EE",X"22",X"F8",X"C8",X"EE",X"22",X"F8",
		X"89",X"EE",X"22",X"F8",X"8F",X"DE",X"77",X"F8",X"8C",X"EE",X"99",X"F8",X"89",X"EE",X"77",X"F8",
		X"89",X"EE",X"66",X"F8",X"89",X"EE",X"66",X"F8",X"99",X"E6",X"66",X"F8",X"FF",X"66",X"66",X"FF",
		X"66",X"66",X"66",X"66",X"66",X"6A",X"66",X"66",X"66",X"6F",X"66",X"66",X"86",X"66",X"66",X"66",
		X"77",X"77",X"88",X"F8",X"77",X"88",X"F9",X"F8",X"77",X"AA",X"CC",X"F8",X"77",X"AA",X"CC",X"F8",
		X"77",X"AA",X"CC",X"F8",X"77",X"AA",X"CC",X"F8",X"F7",X"AA",X"CC",X"F8",X"77",X"AA",X"CC",X"F8",
		X"88",X"AA",X"CC",X"FF",X"88",X"AA",X"CC",X"FC",X"8F",X"AA",X"EE",X"F8",X"88",X"AA",X"CC",X"F8",
		X"89",X"AA",X"CC",X"F8",X"89",X"AA",X"CC",X"F8",X"89",X"AA",X"CC",X"F8",X"89",X"AA",X"CC",X"F8",
		X"7F",X"F7",X"F7",X"F7",X"7F",X"F7",X"F7",X"F7",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"77",X"77",X"77",X"77",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"77",X"77",X"77",X"77",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"F7",X"77",X"77",X"7F",X"F7",X"77",X"77",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"77",X"77",X"77",X"77",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"77",X"77",X"77",X"77",X"FF",X"FF",X"FF",X"FF",
		X"F7",X"66",X"FF",X"FF",X"F7",X"66",X"FF",X"FF",X"F7",X"66",X"FF",X"FF",X"F7",X"66",X"FF",X"FF",
		X"F7",X"66",X"FF",X"FF",X"F7",X"66",X"FF",X"FF",X"F7",X"66",X"FF",X"FF",X"FF",X"66",X"FF",X"FF",
		X"F7",X"66",X"FF",X"FF",X"A7",X"76",X"FF",X"FF",X"66",X"66",X"FF",X"FF",X"66",X"66",X"FF",X"FF",
		X"66",X"6E",X"FF",X"FF",X"66",X"6E",X"FF",X"FF",X"66",X"6F",X"FF",X"FF",X"66",X"EF",X"FF",X"FF",
		X"F7",X"9F",X"66",X"FF",X"F7",X"9F",X"66",X"FF",X"F7",X"9F",X"66",X"FF",X"F7",X"9F",X"66",X"FF",
		X"F7",X"9F",X"66",X"FF",X"F7",X"9F",X"66",X"FF",X"F7",X"9F",X"66",X"FF",X"F7",X"9F",X"66",X"FF",
		X"F7",X"9F",X"66",X"FF",X"F7",X"9F",X"66",X"FF",X"F7",X"9F",X"6D",X"FF",X"F7",X"9F",X"6D",X"FF",
		X"F7",X"F6",X"6F",X"FF",X"F7",X"F6",X"DF",X"FF",X"F7",X"F6",X"DF",X"FF",X"F7",X"66",X"FF",X"FF",
		X"44",X"44",X"44",X"44",X"C4",X"44",X"44",X"44",X"4C",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"44",X"C4",X"44",X"44",X"CC",X"CC",X"CC",X"CC",X"99",X"99",X"99",X"99",X"88",X"88",X"88",X"8F",
		X"88",X"88",X"88",X"8F",X"88",X"88",X"88",X"8F",X"88",X"88",X"88",X"8F",X"FF",X"FF",X"FF",X"FF",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"FF",X"FF",X"FF",X"FF",X"77",X"77",X"77",X"77",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"44",X"44",X"44",X"CC",X"44",X"44",X"44",X"CC",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"C4",X"44",
		X"44",X"44",X"4C",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"C4",X"44",X"44",X"44",X"44",
		X"9F",X"22",X"22",X"F7",X"FF",X"22",X"22",X"F7",X"77",X"22",X"22",X"F7",X"77",X"22",X"2C",X"F7",
		X"79",X"2C",X"CC",X"F9",X"7F",X"EE",X"EE",X"FF",X"7F",X"97",X"77",X"99",X"7F",X"77",X"77",X"77",
		X"7F",X"22",X"22",X"FF",X"77",X"22",X"22",X"F7",X"77",X"22",X"22",X"F7",X"77",X"22",X"22",X"F7",
		X"99",X"E2",X"22",X"F7",X"FF",X"E2",X"22",X"F7",X"7F",X"22",X"22",X"F7",X"7F",X"22",X"22",X"F7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FD",X"FF",X"FF",
		X"FD",X"FF",X"DF",X"EE",X"FF",X"FA",X"DD",X"AA",X"AF",X"FE",X"AE",X"EE",X"AF",X"FE",X"AE",X"EF",
		X"AF",X"FE",X"AE",X"EF",X"AF",X"FE",X"AE",X"EF",X"FF",X"FE",X"AE",X"EF",X"FF",X"FE",X"AE",X"EF",
		X"EA",X"FF",X"AE",X"EF",X"FA",X"FF",X"FE",X"EF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"2C",X"EC",X"AA",X"66",X"88",X"E2",X"9F",X"99",X"88",X"E2",X"9F",X"99",X"88",X"EC",X"9F",
		X"99",X"88",X"EC",X"9F",X"99",X"88",X"EC",X"9F",X"99",X"88",X"EC",X"9F",X"FF",X"AA",X"EC",X"AA",
		X"66",X"99",X"E2",X"66",X"99",X"88",X"EC",X"88",X"99",X"88",X"EC",X"88",X"99",X"88",X"E2",X"88",
		X"99",X"88",X"ED",X"88",X"99",X"88",X"AA",X"88",X"88",X"77",X"CC",X"77",X"66",X"66",X"66",X"66",
		X"FE",X"FE",X"EE",X"AD",X"FF",X"AA",X"EE",X"AE",X"F6",X"FF",X"FF",X"AE",X"F6",X"6F",X"AE",X"FF",
		X"F6",X"6C",X"AE",X"FA",X"F6",X"6F",X"AF",X"FA",X"FC",X"9C",X"FF",X"FF",X"F9",X"8F",X"FF",X"FF",
		X"E8",X"AA",X"EA",X"AA",X"EA",X"AA",X"AA",X"2A",X"EA",X"AA",X"AA",X"CC",X"AA",X"AA",X"2E",X"CC",
		X"AA",X"AA",X"AC",X"CC",X"2A",X"AA",X"2A",X"CC",X"EE",X"EA",X"E2",X"CC",X"66",X"66",X"66",X"66",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"AA",X"FF",X"FF",X"FF",X"AF",X"FF",X"FF",X"FF",X"AE",X"FF",X"FF",X"FF",X"AE",X"FE",X"FF",
		X"FF",X"AE",X"FA",X"AA",X"FF",X"AF",X"FF",X"AA",X"FF",X"AE",X"FF",X"DA",X"FF",X"AE",X"FA",X"DE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"8F",X"FF",X"FF",X"FE",
		X"87",X"AA",X"FF",X"FE",X"87",X"7A",X"FF",X"FE",X"87",X"77",X"FF",X"EE",X"FF",X"FF",X"FF",X"FE",
		X"FA",X"CC",X"CC",X"AC",X"FA",X"CC",X"CC",X"AC",X"FA",X"C2",X"22",X"A2",X"FA",X"C2",X"22",X"A2",
		X"FA",X"C2",X"22",X"A2",X"FA",X"C2",X"22",X"A2",X"FA",X"C2",X"22",X"A2",X"FA",X"C2",X"CC",X"A2",
		X"FA",X"C2",X"CC",X"A2",X"FA",X"C2",X"22",X"A7",X"99",X"99",X"99",X"97",X"F7",X"77",X"77",X"97",
		X"99",X"99",X"99",X"97",X"F7",X"77",X"77",X"97",X"F7",X"77",X"77",X"97",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"CC",X"CC",X"66",X"66",X"CC",X"CC",X"66",X"66",X"CC",X"CC",
		X"66",X"66",X"EE",X"EE",X"EE",X"EE",X"FF",X"FE",X"EE",X"EE",X"FF",X"FF",X"FF",X"FF",X"EE",X"EE",
		X"F9",X"FF",X"FF",X"F9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D5",X"FF",X"FF",X"33",X"DD",X"99",
		X"FF",X"54",X"5D",X"FF",X"FF",X"DD",X"3A",X"FF",X"FF",X"DD",X"3A",X"FF",X"FF",X"5D",X"FF",X"FF",
		X"66",X"66",X"66",X"66",X"66",X"66",X"CC",X"CC",X"66",X"66",X"CC",X"CC",X"66",X"66",X"CC",X"CC",
		X"66",X"66",X"EE",X"EE",X"EE",X"55",X"FF",X"FE",X"EE",X"EE",X"FF",X"FF",X"FF",X"55",X"EE",X"EE",
		X"FC",X"EE",X"FF",X"F9",X"FF",X"EE",X"FF",X"FF",X"FF",X"55",X"BF",X"FF",X"FF",X"EE",X"DB",X"96",
		X"FF",X"55",X"EB",X"FF",X"FF",X"BA",X"BA",X"FF",X"FF",X"AB",X"AE",X"FF",X"FF",X"FA",X"FF",X"FF",
		X"66",X"66",X"DD",X"66",X"66",X"5D",X"DD",X"CC",X"66",X"DD",X"D3",X"CC",X"66",X"DD",X"D5",X"CC",
		X"66",X"F5",X"FE",X"EE",X"EE",X"EF",X"FF",X"FE",X"EE",X"EE",X"FF",X"FF",X"FF",X"FF",X"EE",X"EE",
		X"FF",X"29",X"FB",X"F9",X"FF",X"77",X"99",X"FF",X"FF",X"97",X"79",X"FF",X"FF",X"76",X"9F",X"96",
		X"FF",X"76",X"7A",X"FF",X"FF",X"76",X"7A",X"FF",X"FF",X"77",X"7A",X"FF",X"FF",X"F7",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"CC",X"CC",X"CC",X"CC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"CC",X"CC",X"CC",X"CC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"EE",X"FF",X"FF",X"FF",X"EF",X"FF",X"FF",X"EE",X"FF",X"FF",X"FF",X"EE",X"EE",X"EE",
		X"EE",X"DD",X"DD",X"DD",X"DD",X"DE",X"DD",X"DD",X"DD",X"D6",X"DD",X"DD",X"DD",X"DE",X"DD",X"DD",
		X"AD",X"AA",X"DA",X"DD",X"AD",X"AA",X"AA",X"DD",X"AD",X"AA",X"FF",X"AA",X"AD",X"AA",X"FF",X"FF",
		X"AA",X"AA",X"FF",X"FF",X"FF",X"AA",X"FA",X"FF",X"FF",X"AA",X"FA",X"FF",X"FF",X"FA",X"FF",X"FF",
		X"FF",X"FA",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"DD",X"DD",X"7C",X"77",X"DD",X"D7",X"7C",X"77",X"DD",X"D7",X"CC",X"77",X"AA",X"F7",X"CC",X"77",
		X"A7",X"C7",X"CC",X"77",X"A7",X"C7",X"C7",X"77",X"A7",X"C7",X"C7",X"77",X"A7",X"C7",X"C7",X"77",
		X"77",X"C7",X"C7",X"77",X"77",X"C7",X"C7",X"77",X"7F",X"C7",X"C7",X"77",X"7F",X"C7",X"C7",X"77",
		X"7F",X"C7",X"C7",X"77",X"7F",X"C7",X"C7",X"77",X"7F",X"C7",X"C7",X"77",X"7F",X"C7",X"C7",X"77",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FE",X"EF",
		X"FF",X"FF",X"EF",X"FE",X"FF",X"FE",X"EE",X"ED",X"FF",X"EF",X"DD",X"ED",X"FE",X"EE",X"DD",X"DD",
		X"DD",X"EE",X"FF",X"DD",X"DD",X"DD",X"FF",X"DD",X"DD",X"DD",X"FA",X"DD",X"DD",X"DD",X"DA",X"DD",
		X"DD",X"DD",X"DA",X"DD",X"DD",X"AA",X"DA",X"DD",X"DD",X"FF",X"DA",X"DD",X"DD",X"FF",X"DA",X"DD",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"87",X"FF",X"FF",X"FF",X"77",
		X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"8F",X"77",X"FF",X"FF",X"77",X"77",
		X"FF",X"EE",X"7C",X"77",X"FF",X"EF",X"7C",X"77",X"FF",X"ED",X"7C",X"77",X"EE",X"DD",X"7C",X"77",
		X"77",X"FC",X"C7",X"7C",X"77",X"F7",X"C7",X"7C",X"77",X"F7",X"C7",X"7C",X"77",X"F7",X"C7",X"7C",
		X"77",X"F7",X"C7",X"7C",X"77",X"F7",X"C7",X"7C",X"77",X"F7",X"CC",X"7C",X"77",X"F7",X"C7",X"7C",
		X"77",X"F8",X"C7",X"7C",X"77",X"78",X"C7",X"7C",X"C7",X"78",X"77",X"77",X"C7",X"78",X"77",X"77",
		X"AA",X"78",X"77",X"77",X"AA",X"AA",X"77",X"77",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"11",X"11",X"11",X"1F",X"FF",X"FF",X"FF",X"F1",X"FB",X"BB",X"FB",X"FF",X"FB",X"BF",X"FB",X"FF",
		X"FB",X"BF",X"FB",X"FF",X"FF",X"BF",X"FB",X"FF",X"FF",X"FF",X"FF",X"F1",X"FF",X"1F",X"11",X"18",
		X"FF",X"1F",X"F8",X"88",X"FF",X"FF",X"88",X"88",X"FF",X"FF",X"88",X"88",X"FF",X"FF",X"88",X"88",
		X"FF",X"FF",X"88",X"87",X"FF",X"FF",X"88",X"77",X"FF",X"11",X"99",X"99",X"77",X"99",X"99",X"99",
		X"88",X"11",X"11",X"11",X"88",X"FF",X"FF",X"FF",X"99",X"FF",X"BB",X"BB",X"99",X"FB",X"FF",X"FB",
		X"99",X"FB",X"FF",X"FB",X"99",X"FF",X"BB",X"FB",X"99",X"FF",X"FF",X"FF",X"99",X"11",X"11",X"11",
		X"99",X"FF",X"FF",X"FF",X"99",X"88",X"88",X"FF",X"99",X"88",X"88",X"11",X"99",X"88",X"88",X"FF",
		X"99",X"88",X"87",X"FF",X"99",X"88",X"77",X"FF",X"99",X"99",X"77",X"11",X"99",X"99",X"77",X"88",
		X"66",X"22",X"22",X"F7",X"FF",X"22",X"22",X"F7",X"77",X"22",X"22",X"F7",X"77",X"22",X"22",X"F7",
		X"77",X"22",X"22",X"F7",X"77",X"22",X"22",X"F7",X"77",X"22",X"22",X"F7",X"66",X"CC",X"CC",X"F7",
		X"66",X"88",X"88",X"F7",X"FF",X"22",X"22",X"F7",X"77",X"22",X"22",X"F7",X"77",X"22",X"22",X"F7",
		X"77",X"22",X"22",X"F7",X"77",X"22",X"22",X"F7",X"77",X"22",X"22",X"F7",X"66",X"22",X"22",X"F7",
		X"97",X"7F",X"99",X"7F",X"97",X"7F",X"99",X"7F",X"97",X"7F",X"99",X"7F",X"2A",X"A2",X"AA",X"A2",
		X"22",X"22",X"2E",X"22",X"EE",X"EE",X"EE",X"EE",X"1E",X"E1",X"E1",X"EE",X"EE",X"E1",X"11",X"EE",
		X"1E",X"E1",X"E1",X"EE",X"1E",X"E1",X"E1",X"EE",X"EE",X"EE",X"E1",X"EE",X"3E",X"EE",X"11",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"AA",X"3A",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"77",X"77",X"77",X"77",
		X"FF",X"F7",X"99",X"FF",X"FF",X"97",X"59",X"9F",X"F9",X"57",X"59",X"99",X"F5",X"57",X"59",X"95",
		X"F5",X"57",X"59",X"95",X"F5",X"57",X"59",X"95",X"F5",X"57",X"99",X"95",X"F7",X"77",X"99",X"99",
		X"F7",X"77",X"59",X"99",X"F7",X"57",X"59",X"99",X"F5",X"57",X"59",X"95",X"F5",X"57",X"59",X"95",
		X"F5",X"57",X"59",X"95",X"F5",X"57",X"59",X"95",X"F5",X"57",X"99",X"85",X"F7",X"77",X"99",X"89",
		X"2A",X"CA",X"2A",X"2A",X"2A",X"CA",X"2A",X"2A",X"2A",X"CA",X"CA",X"CA",X"2A",X"CA",X"CA",X"CA",
		X"2A",X"CA",X"CA",X"CA",X"2A",X"CA",X"CA",X"CA",X"2A",X"CA",X"CA",X"CA",X"2A",X"CA",X"CA",X"CA",
		X"2A",X"CA",X"CA",X"CA",X"7A",X"CA",X"CA",X"CA",X"7A",X"CA",X"2A",X"2A",X"FA",X"2A",X"2A",X"2A",
		X"CA",X"2A",X"2A",X"2A",X"CA",X"CA",X"CA",X"CA",X"67",X"77",X"77",X"77",X"66",X"66",X"66",X"66",
		X"77",X"FA",X"88",X"28",X"77",X"FA",X"88",X"28",X"77",X"FA",X"88",X"28",X"77",X"FA",X"88",X"28",
		X"77",X"FA",X"88",X"28",X"77",X"FF",X"89",X"29",X"77",X"FF",X"89",X"29",X"77",X"FF",X"99",X"28",
		X"77",X"FF",X"99",X"28",X"77",X"FF",X"99",X"78",X"77",X"FF",X"99",X"78",X"77",X"6F",X"99",X"C8",
		X"77",X"FF",X"98",X"C8",X"76",X"FF",X"98",X"C8",X"66",X"FF",X"77",X"67",X"FF",X"FF",X"66",X"66",
		X"77",X"FF",X"77",X"77",X"77",X"FF",X"99",X"99",X"77",X"FF",X"88",X"8F",X"77",X"FF",X"77",X"CA",
		X"77",X"FF",X"77",X"2A",X"77",X"FF",X"77",X"2A",X"77",X"FF",X"77",X"2A",X"77",X"FF",X"88",X"88",
		X"77",X"EF",X"99",X"F9",X"77",X"DE",X"88",X"88",X"77",X"DD",X"77",X"C7",X"77",X"DD",X"77",X"C7",
		X"77",X"AA",X"77",X"28",X"77",X"FA",X"78",X"28",X"77",X"FA",X"88",X"28",X"77",X"FA",X"88",X"28",
		X"FF",X"77",X"77",X"77",X"99",X"99",X"99",X"99",X"FF",X"88",X"88",X"87",X"99",X"99",X"99",X"99",
		X"FF",X"88",X"88",X"87",X"99",X"99",X"99",X"99",X"FF",X"88",X"88",X"88",X"99",X"99",X"99",X"FF",
		X"99",X"99",X"99",X"77",X"FF",X"88",X"88",X"77",X"FF",X"FF",X"FF",X"77",X"77",X"77",X"77",X"77",
		X"88",X"88",X"88",X"88",X"99",X"99",X"99",X"99",X"88",X"88",X"88",X"88",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"8F",X"A8",X"FF",X"7F",X"8F",X"8F",X"FF",X"7F",X"8F",X"8F",X"FF",X"7F",X"8F",X"8F",X"FF",
		X"7F",X"8F",X"8F",X"FF",X"7F",X"8F",X"8F",X"FF",X"7F",X"8F",X"8F",X"FF",X"7F",X"8A",X"8F",X"FF",
		X"7F",X"8A",X"8F",X"FF",X"7F",X"AA",X"8F",X"FF",X"7F",X"AA",X"8F",X"FF",X"7F",X"A8",X"8F",X"FF",
		X"7F",X"AF",X"8F",X"FF",X"7F",X"8F",X"8F",X"FF",X"7F",X"8F",X"8F",X"FF",X"7F",X"8F",X"8F",X"FF",
		X"F8",X"77",X"AA",X"AA",X"F9",X"77",X"CC",X"CC",X"F9",X"77",X"CC",X"CC",X"F9",X"77",X"22",X"22",
		X"F9",X"77",X"22",X"22",X"F9",X"77",X"22",X"22",X"F9",X"77",X"A2",X"A2",X"F9",X"77",X"22",X"22",
		X"F9",X"77",X"22",X"22",X"F9",X"77",X"22",X"22",X"F9",X"77",X"22",X"22",X"F9",X"77",X"DD",X"AA",
		X"F9",X"77",X"CC",X"CC",X"F9",X"7C",X"CC",X"CC",X"F8",X"CC",X"CC",X"CC",X"66",X"66",X"66",X"66",
		X"77",X"8F",X"AC",X"FF",X"77",X"8F",X"AC",X"FF",X"77",X"8F",X"AC",X"FF",X"EE",X"8F",X"AC",X"FF",
		X"EE",X"8F",X"AC",X"FF",X"F7",X"8F",X"AC",X"FF",X"F7",X"8F",X"AC",X"8F",X"F7",X"8F",X"AC",X"FF",
		X"F7",X"8F",X"A2",X"FF",X"F7",X"9F",X"AA",X"FF",X"F7",X"9F",X"99",X"FF",X"F7",X"9F",X"77",X"FF",
		X"F7",X"9F",X"DE",X"FF",X"F7",X"9D",X"DD",X"FF",X"F7",X"DD",X"DD",X"FF",X"F7",X"DD",X"DD",X"FF",
		X"FF",X"22",X"FF",X"72",X"FE",X"22",X"EE",X"72",X"F7",X"77",X"77",X"77",X"F7",X"22",X"77",X"72",
		X"F7",X"22",X"88",X"72",X"F7",X"77",X"88",X"77",X"F7",X"22",X"88",X"72",X"F8",X"22",X"88",X"72",
		X"F8",X"77",X"99",X"77",X"F8",X"22",X"99",X"72",X"F9",X"22",X"99",X"7C",X"F9",X"77",X"99",X"77",
		X"F9",X"22",X"99",X"7C",X"F9",X"CC",X"99",X"7C",X"F9",X"77",X"99",X"77",X"F9",X"CC",X"99",X"7C",
		X"F8",X"88",X"88",X"88",X"8A",X"CC",X"AF",X"AA",X"7A",X"CC",X"AF",X"CC",X"7A",X"CC",X"A7",X"CC",
		X"7A",X"22",X"A7",X"2C",X"7A",X"22",X"A7",X"2C",X"7A",X"22",X"A7",X"2C",X"7A",X"22",X"A7",X"2C",
		X"7A",X"22",X"A7",X"2C",X"7A",X"22",X"A7",X"2C",X"7A",X"22",X"A7",X"2C",X"7A",X"CC",X"A7",X"2C",
		X"7A",X"22",X"AC",X"CC",X"7A",X"FF",X"CC",X"CC",X"CA",X"CC",X"CC",X"AA",X"66",X"66",X"66",X"66",
		X"44",X"77",X"07",X"F7",X"44",X"47",X"F7",X"F7",X"74",X"47",X"00",X"F7",X"74",X"47",X"F7",X"F7",
		X"74",X"77",X"07",X"F7",X"44",X"44",X"F0",X"F7",X"44",X"44",X"00",X"F7",X"77",X"77",X"F7",X"F7",
		X"44",X"44",X"00",X"F7",X"44",X"44",X"F7",X"F7",X"74",X"47",X"00",X"F7",X"74",X"47",X"F7",X"F7",
		X"44",X"47",X"00",X"F7",X"44",X"47",X"F7",X"F7",X"FF",X"FF",X"00",X"FF",X"77",X"77",X"F7",X"F7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"4F",X"F4",X"FF",X"FF",X"FF",X"4F",
		X"FF",X"FF",X"4F",X"44",X"FF",X"FF",X"FF",X"4F",X"FF",X"FF",X"FF",X"4F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",
		X"88",X"88",X"88",X"18",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",
		X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",
		X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",
		X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DD",X"DD",X"DD",
		X"DD",X"D5",X"5D",X"55",X"79",X"AC",X"CA",X"CC",X"79",X"AC",X"CA",X"CC",X"79",X"A5",X"5A",X"55",
		X"79",X"A5",X"5A",X"55",X"79",X"A5",X"5A",X"55",X"79",X"A5",X"5A",X"55",X"79",X"A5",X"CA",X"CC",
		X"79",X"A5",X"CA",X"CC",X"79",X"A5",X"CA",X"CC",X"78",X"88",X"88",X"88",X"77",X"AE",X"EE",X"EE",
		X"7F",X"F7",X"F7",X"F7",X"7F",X"F7",X"F7",X"F7",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"77",X"77",X"77",X"77",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"77",X"77",X"77",X"77",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"F7",X"77",X"77",X"7F",X"F7",X"77",X"77",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"77",X"77",X"77",X"77",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"33",X"33",X"33",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"77",X"77",X"77",X"77",X"FF",X"FF",X"FF",X"FF",
		X"66",X"22",X"22",X"F7",X"FF",X"22",X"22",X"F7",X"70",X"CC",X"00",X"47",X"70",X"C2",X"CC",X"F4",
		X"70",X"C2",X"22",X"F4",X"70",X"CC",X"22",X"F4",X"70",X"00",X"22",X"F4",X"66",X"CC",X"CC",X"F4",
		X"66",X"88",X"88",X"F4",X"44",X"44",X"44",X"47",X"77",X"CC",X"CC",X"F7",X"77",X"2C",X"C2",X"F7",
		X"44",X"2C",X"C2",X"F7",X"77",X"CC",X"CC",X"47",X"44",X"44",X"44",X"F7",X"66",X"CC",X"CC",X"F7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"4F",X"44",X"44",X"FF",X"FF",X"4F",X"FF",X"FF",
		X"FF",X"44",X"44",X"FF",X"FF",X"4F",X"F4",X"FF",X"FF",X"44",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"11",X"11",X"FF",X"FF",X"1F",X"FF",X"FF",X"FF",X"1F",X"1F",X"FF",X"FF",X"1F",X"F1",X"FF",X"FF",
		X"11",X"18",X"88",X"88",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",
		X"FF",X"FC",X"FF",X"FF",X"99",X"9C",X"99",X"FF",X"79",X"99",X"99",X"FF",X"99",X"99",X"98",X"FF",
		X"98",X"98",X"99",X"FF",X"99",X"99",X"88",X"FF",X"FF",X"99",X"FC",X"FF",X"8C",X"FF",X"FC",X"FF",
		X"9C",X"CF",X"FC",X"FF",X"99",X"CF",X"FC",X"FF",X"99",X"FC",X"FC",X"FF",X"99",X"98",X"FC",X"7F",
		X"99",X"9F",X"F2",X"7F",X"99",X"8F",X"F2",X"FF",X"99",X"7F",X"FF",X"FF",X"99",X"7F",X"99",X"FF",
		X"78",X"CC",X"CC",X"88",X"78",X"CC",X"CC",X"88",X"78",X"22",X"22",X"88",X"79",X"2C",X"2C",X"99",
		X"79",X"CC",X"2C",X"99",X"79",X"CC",X"22",X"99",X"79",X"CC",X"2C",X"99",X"79",X"CC",X"2C",X"99",
		X"79",X"CC",X"2C",X"99",X"79",X"CC",X"2C",X"99",X"79",X"CC",X"CC",X"99",X"79",X"CC",X"2C",X"99",
		X"79",X"CC",X"CC",X"99",X"79",X"99",X"99",X"99",X"79",X"77",X"77",X"99",X"66",X"66",X"66",X"66",
		X"77",X"55",X"77",X"55",X"77",X"55",X"77",X"55",X"77",X"5F",X"77",X"55",X"77",X"5F",X"F5",X"55",
		X"77",X"5F",X"F5",X"55",X"77",X"5F",X"F5",X"55",X"77",X"5F",X"F5",X"55",X"77",X"5F",X"FF",X"FF",
		X"77",X"F7",X"BB",X"7B",X"77",X"77",X"BB",X"BB",X"77",X"77",X"3F",X"33",X"77",X"77",X"33",X"33",
		X"77",X"77",X"33",X"33",X"77",X"77",X"4F",X"44",X"77",X"77",X"44",X"44",X"77",X"77",X"44",X"44",
		X"77",X"77",X"77",X"77",X"75",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"75",X"55",X"5F",X"75",
		X"75",X"FF",X"55",X"5F",X"75",X"55",X"55",X"5F",X"55",X"55",X"55",X"5F",X"FF",X"FF",X"FF",X"FF",
		X"7B",X"BF",X"BB",X"55",X"7B",X"BF",X"BB",X"5F",X"7F",X"F7",X"33",X"5F",X"77",X"77",X"33",X"77",
		X"77",X"77",X"33",X"77",X"77",X"77",X"44",X"77",X"77",X"77",X"44",X"77",X"77",X"77",X"44",X"77",
		X"FF",X"FF",X"FF",X"FF",X"99",X"99",X"9F",X"99",X"77",X"FF",X"F9",X"97",X"88",X"99",X"F9",X"99",
		X"88",X"99",X"99",X"99",X"99",X"89",X"98",X"77",X"79",X"89",X"99",X"88",X"87",X"99",X"99",X"88",
		X"87",X"99",X"99",X"88",X"99",X"99",X"77",X"99",X"99",X"7F",X"99",X"99",X"FF",X"88",X"99",X"9F",
		X"99",X"98",X"99",X"99",X"99",X"99",X"99",X"99",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"FF",X"F6",X"66",X"66",X"FF",X"66",X"66",X"66",X"FF",X"66",X"66",X"66",X"FF",X"88",X"88",X"88",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"88",X"88",X"88",X"88",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F7",X"78",X"99",X"89",X"F7",X"78",X"99",X"89",X"F7",X"78",X"99",X"89",X"FA",X"A2",X"AA",X"A2",
		X"FE",X"22",X"2E",X"E2",X"FE",X"EE",X"EE",X"EE",X"FE",X"EE",X"1E",X"EE",X"FE",X"EE",X"E1",X"EE",
		X"FE",X"EE",X"1E",X"EE",X"FE",X"EE",X"EE",X"11",X"FE",X"EE",X"EE",X"EE",X"FE",X"EE",X"EE",X"33",
		X"FE",X"EE",X"EE",X"3E",X"FA",X"AA",X"AA",X"33",X"FF",X"FF",X"FF",X"FF",X"F7",X"77",X"77",X"77",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"88",X"88",X"88",X"88",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F7",X"77",X"99",X"89",X"F7",X"77",X"99",X"89",X"F7",X"77",X"99",X"89",X"F7",X"77",X"99",X"89",
		X"F7",X"77",X"99",X"89",X"F7",X"77",X"99",X"89",X"F7",X"77",X"99",X"89",X"F7",X"77",X"99",X"89",
		X"F7",X"77",X"99",X"89",X"FA",X"77",X"99",X"AE",X"F7",X"AA",X"DD",X"89",X"F7",X"77",X"77",X"89",
		X"F7",X"87",X"77",X"89",X"F7",X"88",X"78",X"89",X"C7",X"CC",X"CC",X"89",X"66",X"66",X"66",X"66",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",
		X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",
		X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",
		X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"99",X"FF",X"FF",X"FF",X"55",X"FF",X"FF",X"FF",X"55",
		X"FF",X"FF",X"FF",X"55",X"FF",X"FF",X"FF",X"99",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"D7",X"EA",X"7E",X"FF",X"D7",X"7A",X"7E",X"FF",X"D7",X"F7",X"7F",X"FA",X"F7",X"FA",X"7F",X"FA",
		X"C7",X"FA",X"7F",X"FA",X"99",X"99",X"99",X"FF",X"88",X"88",X"89",X"FF",X"99",X"99",X"88",X"6F",
		X"88",X"88",X"98",X"99",X"88",X"88",X"98",X"88",X"77",X"78",X"98",X"88",X"77",X"77",X"98",X"88",
		X"77",X"77",X"98",X"88",X"77",X"77",X"98",X"78",X"77",X"77",X"97",X"77",X"FF",X"FF",X"FA",X"FF",
		X"99",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"90",X"F0",X"FF",X"F0",X"70",X"F0",X"0F",X"0F",
		X"99",X"F0",X"0F",X"09",X"77",X"90",X"0F",X"07",X"99",X"70",X"FF",X"70",X"99",X"97",X"FF",X"97",
		X"77",X"39",X"33",X"39",X"77",X"97",X"37",X"38",X"77",X"39",X"33",X"79",X"77",X"99",X"99",X"99",
		X"88",X"FF",X"FF",X"FF",X"99",X"99",X"99",X"99",X"88",X"88",X"88",X"88",X"FF",X"FF",X"FF",X"FF",
		X"88",X"8F",X"88",X"88",X"8F",X"F8",X"2C",X"CA",X"F8",X"88",X"CC",X"A8",X"F7",X"77",X"FA",X"F7",
		X"F7",X"77",X"CA",X"A7",X"F7",X"77",X"CA",X"A7",X"F7",X"77",X"CA",X"A7",X"F7",X"77",X"CA",X"A7",
		X"F7",X"77",X"CA",X"A7",X"F7",X"77",X"2A",X"A7",X"F7",X"77",X"2A",X"A7",X"F7",X"77",X"2A",X"A7",
		X"F7",X"77",X"2A",X"A7",X"F7",X"77",X"2A",X"A7",X"F7",X"77",X"2A",X"A7",X"F7",X"77",X"2A",X"A7",
		X"88",X"88",X"88",X"88",X"A8",X"88",X"8A",X"22",X"88",X"88",X"AA",X"CC",X"77",X"77",X"A0",X"FF",
		X"77",X"77",X"AC",X"CC",X"77",X"77",X"AC",X"CC",X"77",X"77",X"EC",X"22",X"77",X"77",X"EC",X"22",
		X"77",X"77",X"EC",X"22",X"77",X"77",X"EC",X"22",X"77",X"77",X"EC",X"22",X"77",X"77",X"EC",X"22",
		X"77",X"77",X"EC",X"22",X"77",X"77",X"EC",X"22",X"77",X"77",X"E2",X"22",X"77",X"77",X"A2",X"22",
		X"C7",X"87",X"66",X"9F",X"C8",X"88",X"66",X"9F",X"CC",X"88",X"67",X"9F",X"88",X"88",X"66",X"FF",
		X"88",X"88",X"76",X"7F",X"88",X"88",X"67",X"9F",X"88",X"88",X"66",X"9F",X"88",X"88",X"66",X"9F",
		X"88",X"88",X"66",X"9F",X"88",X"88",X"F6",X"8F",X"88",X"88",X"C6",X"8F",X"FF",X"88",X"66",X"8F",
		X"AA",X"77",X"66",X"8F",X"CA",X"FF",X"66",X"8F",X"CC",X"AA",X"66",X"8F",X"CA",X"AA",X"66",X"7F",
		X"AA",X"AA",X"A6",X"AA",X"77",X"77",X"66",X"77",X"77",X"7A",X"66",X"7A",X"7A",X"AF",X"66",X"AF",
		X"7A",X"AF",X"66",X"AF",X"7A",X"AF",X"66",X"AC",X"7A",X"AF",X"66",X"AC",X"7A",X"AF",X"66",X"AC",
		X"CC",X"AF",X"6F",X"A2",X"7C",X"AF",X"66",X"A2",X"7C",X"AF",X"66",X"A2",X"7C",X"AF",X"88",X"A2",
		X"FC",X"ED",X"66",X"A2",X"CC",X"88",X"66",X"EE",X"FF",X"77",X"66",X"77",X"77",X"87",X"66",X"99",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",X"6F",X"77",X"FF",X"AA",X"7F",X"77",
		X"FF",X"88",X"FC",X"77",X"AA",X"88",X"C9",X"77",X"88",X"88",X"77",X"7F",X"88",X"8A",X"77",X"F8",
		X"88",X"8A",X"77",X"88",X"88",X"7A",X"F7",X"F8",X"88",X"7A",X"6F",X"F8",X"87",X"7A",X"86",X"F8",
		X"77",X"7A",X"86",X"F8",X"76",X"7A",X"86",X"F8",X"17",X"6F",X"81",X"F8",X"77",X"77",X"66",X"77",
		X"CC",X"FF",X"EF",X"DD",X"11",X"11",X"F1",X"11",X"F1",X"E1",X"81",X"18",X"91",X"11",X"F1",X"F8",
		X"91",X"1F",X"F1",X"F8",X"91",X"F1",X"11",X"F6",X"98",X"88",X"88",X"86",X"98",X"17",X"1F",X"F1",
		X"FF",X"F1",X"1F",X"F1",X"FF",X"F1",X"1F",X"1F",X"FF",X"F1",X"1F",X"1F",X"AA",X"17",X"1F",X"1F",
		X"AC",X"88",X"88",X"AF",X"CC",X"AC",X"CF",X"77",X"CC",X"9C",X"CF",X"77",X"CC",X"9C",X"FC",X"77",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",
		X"FF",X"FF",X"FC",X"CC",X"FF",X"FF",X"FC",X"CF",X"FF",X"FF",X"FC",X"CF",X"FF",X"FF",X"77",X"77",
		X"DD",X"AA",X"FF",X"FF",X"DD",X"FF",X"AF",X"FF",X"FD",X"FF",X"FD",X"FA",X"FF",X"FF",X"FD",X"FA",
		X"FF",X"FF",X"FF",X"D6",X"FF",X"FF",X"FF",X"69",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",
		X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"66",X"67",X"FF",X"AA",X"76",X"79",X"FC",X"AA",X"77",X"7C",
		X"AA",X"CC",X"77",X"7C",X"AC",X"C7",X"97",X"7F",X"CC",X"FF",X"FF",X"FF",X"CC",X"CC",X"CC",X"CC",
		X"FF",X"FF",X"AA",X"AA",X"FF",X"FF",X"FF",X"CC",X"FF",X"FF",X"FF",X"CF",X"FF",X"FF",X"FF",X"CC",
		X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",
		X"FF",X"FF",X"FF",X"CF",X"FF",X"7F",X"FF",X"CF",X"FF",X"9F",X"FF",X"CF",X"FF",X"99",X"FF",X"CF",
		X"FF",X"99",X"FF",X"CC",X"DF",X"2F",X"FF",X"FC",X"DD",X"FF",X"FF",X"FC",X"DD",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"66",X"AA",X"AA",X"AA",X"AA",X"AC",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AE",X"AA",X"CA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EE",X"AA",X"AA",X"AA",X"ED",X"AA",X"AA",
		X"AA",X"FE",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AE",X"AA",X"AA",
		X"AA",X"EE",X"AD",X"AA",X"AA",X"AA",X"AA",X"AA",X"CC",X"66",X"CC",X"CC",X"CF",X"6C",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"AC",X"CC",X"CC",X"CC",X"AA",X"CC",X"CC",X"CC",
		X"AA",X"CC",X"CC",X"CC",X"AA",X"CC",X"CC",X"CC",X"CA",X"CC",X"8C",X"CC",X"CA",X"AA",X"CC",X"CA",
		X"FC",X"AE",X"CC",X"AA",X"FC",X"AA",X"AA",X"AA",X"FF",X"AA",X"CA",X"AA",X"FF",X"AA",X"AA",X"EE",
		X"FF",X"AA",X"AA",X"FE",X"FF",X"FF",X"AA",X"AA",X"FF",X"FC",X"CC",X"CC",X"FF",X"CC",X"CC",X"C6",
		X"CC",X"9C",X"EC",X"77",X"CC",X"9C",X"CC",X"77",X"FF",X"9F",X"FF",X"77",X"FF",X"7C",X"CC",X"CC",
		X"AA",X"CC",X"CC",X"AA",X"AA",X"CC",X"CC",X"AA",X"AA",X"AA",X"CC",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"DE",X"AA",X"AA",X"AA",X"AE",X"AA",X"AA",X"DA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AD",X"AA",X"AA",X"AA",X"FF",X"CC",X"CE",X"66",X"FC",X"CC",X"CC",X"66",
		X"FF",X"77",X"FF",X"FF",X"FF",X"70",X"77",X"1F",X"FF",X"70",X"70",X"FF",X"FF",X"70",X"70",X"1F",
		X"FF",X"70",X"70",X"1F",X"FF",X"70",X"70",X"FF",X"FF",X"70",X"70",X"FF",X"FF",X"70",X"70",X"44",
		X"F8",X"70",X"70",X"F4",X"F8",X"70",X"70",X"F4",X"F8",X"70",X"70",X"F4",X"F8",X"70",X"70",X"84",
		X"F8",X"70",X"70",X"88",X"F8",X"70",X"70",X"88",X"F8",X"70",X"70",X"88",X"76",X"2F",X"2F",X"66",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"96",X"FF",X"FF",X"A7",X"67",X"FF",X"AA",X"77",X"67",
		X"FF",X"88",X"77",X"97",X"AA",X"88",X"77",X"77",X"88",X"88",X"77",X"7F",X"88",X"8A",X"77",X"F8",
		X"88",X"8A",X"77",X"88",X"88",X"7A",X"F7",X"F8",X"88",X"7A",X"6F",X"F8",X"87",X"7A",X"86",X"F8",
		X"77",X"7A",X"86",X"F8",X"76",X"7A",X"86",X"F8",X"17",X"6F",X"81",X"F8",X"77",X"77",X"66",X"77",
		X"AA",X"FF",X"FC",X"AA",X"AA",X"FF",X"FC",X"AA",X"AC",X"FF",X"FF",X"AA",X"AC",X"FF",X"FF",X"CC",
		X"CF",X"FF",X"FF",X"FF",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"DD",X"DD",X"DD",X"AF",X"DD",X"DD",X"AD",X"AF",X"AA",X"AA",X"AD",X"FF",X"FA",X"AF",X"AD",
		X"FF",X"FF",X"FF",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",
		X"FF",X"7F",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"F2",X"7F",X"FF",X"FF",X"FF",X"AA",X"AA",X"AA",
		X"CF",X"FC",X"AA",X"AA",X"AC",X"FF",X"AA",X"AA",X"AA",X"FF",X"AA",X"AA",X"AA",X"FF",X"CA",X"AA",
		X"66",X"66",X"66",X"66",X"66",X"EE",X"66",X"66",X"66",X"66",X"66",X"66",X"88",X"88",X"88",X"88",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"99",X"99",X"9F",X"FF",X"77",X"77",X"8F",X"FF",
		X"88",X"88",X"8F",X"FF",X"88",X"88",X"FF",X"FF",X"88",X"88",X"FF",X"FF",X"88",X"8F",X"FF",X"FF",
		X"88",X"6F",X"CF",X"FF",X"87",X"6F",X"8F",X"FF",X"88",X"FF",X"8F",X"FF",X"88",X"8F",X"8F",X"FF",
		X"F7",X"ED",X"DD",X"FF",X"F7",X"ED",X"DD",X"FF",X"F7",X"EE",X"DD",X"FF",X"F7",X"EE",X"DD",X"FF",
		X"F7",X"EE",X"DD",X"FF",X"F7",X"EE",X"DD",X"66",X"F7",X"EE",X"DD",X"66",X"F7",X"EE",X"DD",X"66",
		X"F7",X"EE",X"DD",X"6D",X"F7",X"EE",X"DD",X"6D",X"F7",X"EE",X"DD",X"6F",X"F7",X"EE",X"DD",X"DF",
		X"F7",X"EE",X"DD",X"DF",X"F7",X"9E",X"DD",X"FF",X"F7",X"9F",X"D6",X"FF",X"F7",X"9F",X"66",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",
		X"F7",X"9F",X"DE",X"FF",X"77",X"9D",X"DD",X"FF",X"F9",X"DD",X"DD",X"FF",X"F9",X"DD",X"DD",X"FF",
		X"F7",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"7F",X"77",X"FA",X"FF",X"7F",X"77",X"EA",X"FF",X"78",
		X"77",X"DE",X"ED",X"F9",X"77",X"DA",X"FF",X"F9",X"77",X"EA",X"FF",X"F9",X"77",X"EA",X"FF",X"F9",
		X"77",X"EA",X"FF",X"F9",X"99",X"EA",X"FF",X"FF",X"99",X"EA",X"FF",X"F7",X"99",X"EA",X"FF",X"F8",
		X"99",X"EA",X"FF",X"F8",X"98",X"EA",X"EE",X"F8",X"8F",X"EE",X"AA",X"F8",X"FF",X"F9",X"FF",X"F8",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"88",X"88",X"88",X"88",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"99",X"99",X"FF",X"99",X"77",X"77",
		X"FF",X"77",X"88",X"88",X"FF",X"88",X"88",X"68",X"99",X"FC",X"88",X"88",X"77",X"FA",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"99",X"88",X"99",X"96",X"77",X"99",X"77",
		X"66",X"66",X"66",X"66",X"66",X"66",X"CC",X"CC",X"66",X"66",X"CC",X"CC",X"66",X"66",X"CC",X"CC",
		X"66",X"66",X"EE",X"EE",X"EE",X"EE",X"F1",X"FE",X"EE",X"EE",X"F8",X"FF",X"FF",X"FF",X"EE",X"EE",
		X"F9",X"FF",X"FF",X"F9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DD",X"99",
		X"FF",X"5D",X"DD",X"FF",X"FF",X"DD",X"DD",X"FF",X"FF",X"DD",X"D5",X"FF",X"FF",X"F5",X"FF",X"FF",
		X"66",X"FF",X"FF",X"FF",X"66",X"CF",X"FF",X"FF",X"66",X"FF",X"FF",X"FF",X"66",X"C8",X"FF",X"FF",
		X"66",X"FF",X"FF",X"FF",X"EE",X"FF",X"FF",X"FF",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"88",X"88",X"88",X"88",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"99",X"99",X"99",X"99",X"77",X"77",X"77",X"7C",
		X"88",X"88",X"88",X"8C",X"88",X"88",X"A9",X"FC",X"88",X"8A",X"99",X"8F",X"8F",X"CC",X"98",X"88",
		X"88",X"CC",X"88",X"77",X"88",X"88",X"88",X"78",X"79",X"78",X"89",X"88",X"97",X"99",X"97",X"99",
		X"88",X"8F",X"8F",X"FF",X"E8",X"8F",X"8F",X"FF",X"FE",X"8F",X"8C",X"FF",X"FE",X"8F",X"87",X"FF",
		X"FC",X"8F",X"8C",X"FF",X"CF",X"8F",X"8C",X"FF",X"7F",X"8F",X"89",X"FF",X"7F",X"8F",X"89",X"FF",
		X"7F",X"8F",X"89",X"FF",X"7F",X"CF",X"89",X"FF",X"7F",X"9F",X"89",X"FF",X"7F",X"7F",X"8D",X"FF",
		X"7F",X"7F",X"8A",X"FF",X"7F",X"8F",X"8A",X"FF",X"7F",X"8F",X"AA",X"FF",X"7F",X"8F",X"AF",X"FF",
		X"99",X"55",X"99",X"99",X"77",X"55",X"FF",X"FF",X"77",X"FF",X"5F",X"55",X"77",X"77",X"5F",X"FF",
		X"77",X"55",X"5F",X"55",X"77",X"FF",X"5F",X"FF",X"77",X"55",X"55",X"55",X"77",X"55",X"55",X"55",
		X"77",X"22",X"FF",X"FF",X"77",X"2F",X"F5",X"55",X"77",X"F5",X"5F",X"55",X"77",X"2F",X"F5",X"FF",
		X"77",X"2F",X"F5",X"5F",X"77",X"F5",X"5F",X"5F",X"77",X"5F",X"2F",X"F2",X"77",X"F5",X"F5",X"22",
		X"77",X"8F",X"85",X"55",X"77",X"8F",X"85",X"5F",X"77",X"8F",X"85",X"55",X"EE",X"8F",X"85",X"5F",
		X"EE",X"8F",X"85",X"5F",X"F8",X"8F",X"8F",X"FF",X"F8",X"8F",X"85",X"55",X"F8",X"8F",X"95",X"F5",
		X"F8",X"9F",X"95",X"55",X"F8",X"9F",X"9F",X"FF",X"F8",X"9F",X"9F",X"FF",X"F8",X"9F",X"9F",X"FF",
		X"F8",X"9F",X"DE",X"FF",X"F8",X"9D",X"DD",X"FF",X"F8",X"DD",X"DD",X"FF",X"F7",X"DD",X"DD",X"FF",
		X"F7",X"DD",X"DD",X"FF",X"F7",X"DD",X"DD",X"FF",X"F7",X"DD",X"DD",X"FF",X"F7",X"DD",X"DD",X"FF",
		X"F7",X"DD",X"DD",X"FF",X"F7",X"DD",X"DD",X"FF",X"F7",X"DD",X"DD",X"FF",X"F7",X"DD",X"DD",X"FF",
		X"F7",X"DD",X"DD",X"FF",X"F7",X"DD",X"DD",X"FF",X"F7",X"DD",X"DD",X"FF",X"F7",X"DD",X"DD",X"FF",
		X"F7",X"DD",X"DD",X"FF",X"F7",X"DD",X"DD",X"FF",X"F7",X"DD",X"DD",X"FF",X"F7",X"DD",X"DD",X"FF",
		X"99",X"99",X"99",X"99",X"FF",X"FF",X"FF",X"FF",X"55",X"55",X"55",X"55",X"FF",X"F7",X"F5",X"FF",
		X"F7",X"F2",X"55",X"55",X"FF",X"FF",X"5F",X"FF",X"55",X"55",X"F5",X"FF",X"55",X"55",X"F5",X"FF",
		X"FF",X"FF",X"2F",X"FF",X"55",X"55",X"5F",X"55",X"55",X"55",X"55",X"FF",X"F5",X"FF",X"55",X"5F",
		X"F5",X"55",X"5F",X"5F",X"F5",X"55",X"5F",X"FF",X"55",X"FF",X"5F",X"55",X"55",X"FF",X"5F",X"5F",
		X"F7",X"FF",X"22",X"F7",X"F7",X"CF",X"22",X"F7",X"F7",X"77",X"22",X"F7",X"EE",X"E7",X"2C",X"EE",
		X"EE",X"D7",X"FF",X"AA",X"77",X"D7",X"FF",X"AA",X"77",X"DA",X"AA",X"AF",X"77",X"EE",X"AA",X"FC",
		X"77",X"77",X"7F",X"F7",X"77",X"77",X"F7",X"F7",X"77",X"FF",X"FF",X"F7",X"77",X"AA",X"AA",X"F7",
		X"77",X"FF",X"CC",X"F7",X"77",X"FF",X"CC",X"F7",X"77",X"FF",X"CC",X"F8",X"F7",X"FA",X"22",X"F8");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
