library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity turkey_shoot_graph3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of turkey_shoot_graph3 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"78",X"FF",X"FF",X"FF",X"78",X"FF",X"FF",X"FF",X"78",X"FF",X"FF",X"FF",X"78",X"FF",X"EE",X"FF",
		X"78",X"22",X"22",X"FF",X"78",X"2A",X"2C",X"FF",X"78",X"DE",X"AA",X"FF",X"77",X"AC",X"DD",X"FF",
		X"77",X"A2",X"CC",X"AC",X"77",X"AA",X"EE",X"AC",X"77",X"CA",X"AA",X"CC",X"77",X"7A",X"77",X"7C",
		X"77",X"CC",X"CC",X"CC",X"77",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"66",X"66",X"66",X"66",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"F3",X"F3",X"FF",X"F3",X"F3",X"3F",X"FF",X"F3",X"F3",X"F3",
		X"F3",X"F3",X"F3",X"FF",X"FF",X"3F",X"F3",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",
		X"FF",X"FF",X"F1",X"1F",X"FF",X"FF",X"F1",X"11",X"FF",X"FF",X"F1",X"1F",X"FF",X"FF",X"FF",X"1F",
		X"7F",X"7F",X"77",X"77",X"7F",X"7F",X"77",X"77",X"7F",X"7F",X"77",X"77",X"7F",X"7F",X"77",X"77",
		X"7F",X"7F",X"77",X"77",X"7F",X"7F",X"77",X"77",X"7F",X"7F",X"77",X"77",X"7F",X"7F",X"77",X"77",
		X"7F",X"7F",X"77",X"77",X"7F",X"7F",X"77",X"77",X"7F",X"7F",X"77",X"77",X"7F",X"7F",X"77",X"77",
		X"7F",X"7F",X"77",X"77",X"7F",X"7F",X"77",X"77",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"77",X"77",
		X"7F",X"F7",X"FF",X"FF",X"9C",X"C9",X"FF",X"CF",X"88",X"88",X"FF",X"88",X"5C",X"F5",X"5C",X"5C",
		X"5C",X"5C",X"CC",X"CC",X"5C",X"FC",X"CC",X"CC",X"FC",X"55",X"CC",X"5C",X"88",X"88",X"88",X"88",
		X"99",X"99",X"99",X"99",X"88",X"88",X"88",X"88",X"FC",X"FC",X"CC",X"CC",X"FC",X"FC",X"CC",X"CC",
		X"F2",X"F2",X"22",X"22",X"F2",X"F2",X"22",X"22",X"F2",X"F2",X"22",X"22",X"F2",X"F2",X"22",X"22",
		X"77",X"F7",X"7F",X"77",X"F9",X"99",X"9F",X"99",X"88",X"88",X"FF",X"88",X"72",X"72",X"72",X"72",
		X"72",X"75",X"72",X"72",X"72",X"75",X"72",X"72",X"72",X"75",X"55",X"72",X"F8",X"88",X"FF",X"88",
		X"99",X"99",X"FF",X"99",X"88",X"88",X"FF",X"88",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"72",X"72",X"72",X"72",X"A2",X"A2",X"A2",X"A2",X"A2",X"A2",X"A2",X"A2",X"A2",X"A2",X"A2",X"A2",
		X"FD",X"FF",X"FF",X"DF",X"FF",X"FF",X"FD",X"DD",X"FF",X"FD",X"FF",X"DD",X"FF",X"DD",X"DF",X"DD",
		X"FF",X"DD",X"33",X"DD",X"FF",X"33",X"FF",X"33",X"DD",X"FF",X"11",X"FF",X"EE",X"FF",X"FF",X"1F",
		X"FD",X"1F",X"FF",X"F1",X"DE",X"F1",X"FF",X"FF",X"DD",X"FF",X"11",X"FF",X"DD",X"FF",X"FF",X"FF",
		X"DD",X"FF",X"FF",X"F1",X"EE",X"FF",X"FF",X"1F",X"EE",X"FF",X"33",X"FF",X"EE",X"33",X"EF",X"33",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"D3",X"FF",X"FF",X"F3",X"3F",X"3F",X"FF",X"1F",X"FF",X"3F",X"FF",X"1F",X"F1",X"3F",X"FF",
		X"1F",X"F1",X"3E",X"FF",X"1F",X"FF",X"3D",X"FF",X"1F",X"FF",X"3E",X"FD",X"1F",X"F1",X"3E",X"DD",
		X"1F",X"FF",X"3D",X"DD",X"FF",X"FF",X"3E",X"DD",X"3F",X"F3",X"EE",X"DE",X"D3",X"3D",X"EE",X"EE",
		X"77",X"77",X"77",X"22",X"B1",X"B1",X"B1",X"22",X"22",X"22",X"22",X"22",X"11",X"11",X"22",X"22",
		X"FF",X"FF",X"12",X"22",X"11",X"F2",X"1F",X"F2",X"FF",X"F2",X"1F",X"22",X"11",X"F2",X"1F",X"F2",
		X"FF",X"F2",X"2F",X"F2",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"B1",X"B1",X"B1",X"B1",
		X"77",X"FF",X"FF",X"77",X"77",X"AA",X"AA",X"77",X"99",X"CA",X"CA",X"99",X"99",X"CA",X"CA",X"99",
		X"77",X"77",X"77",X"8F",X"B1",X"B1",X"B1",X"8F",X"22",X"22",X"22",X"BF",X"22",X"12",X"21",X"21",
		X"12",X"F1",X"F1",X"2B",X"2F",X"21",X"21",X"21",X"12",X"21",X"F1",X"2B",X"1F",X"12",X"21",X"21",
		X"2F",X"FF",X"F2",X"2B",X"22",X"22",X"22",X"21",X"22",X"22",X"22",X"BF",X"B1",X"B1",X"B1",X"8F",
		X"FF",X"FF",X"FF",X"9F",X"AA",X"AA",X"FF",X"9F",X"CC",X"CC",X"F7",X"9F",X"CC",X"CC",X"77",X"9F",
		X"7F",X"CC",X"22",X"66",X"7F",X"00",X"CC",X"FF",X"7F",X"0C",X"00",X"07",X"7F",X"0C",X"0C",X"70",
		X"7F",X"0C",X"00",X"70",X"7F",X"0C",X"0C",X"00",X"7F",X"0C",X"00",X"70",X"7F",X"CC",X"CC",X"77",
		X"74",X"44",X"77",X"77",X"74",X"4C",X"24",X"44",X"74",X"4C",X"4C",X"47",X"74",X"4C",X"4C",X"47",
		X"74",X"4C",X"4C",X"44",X"74",X"4C",X"4C",X"47",X"7F",X"4C",X"C4",X"44",X"7F",X"C2",X"2C",X"77",
		X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"07",X"FF",X"FF",X"77",X"07",X"FF",X"FF",X"07",X"07",X"FF",
		X"FF",X"07",X"07",X"FF",X"1F",X"07",X"07",X"FF",X"FF",X"07",X"07",X"FF",X"4F",X"07",X"07",X"8F",
		X"F4",X"07",X"07",X"8F",X"4F",X"07",X"07",X"8F",X"F4",X"07",X"07",X"8F",X"74",X"07",X"07",X"8F",
		X"88",X"07",X"07",X"8F",X"88",X"07",X"07",X"8F",X"EE",X"07",X"07",X"EA",X"66",X"F2",X"F2",X"67",
		X"00",X"FF",X"FF",X"FF",X"F4",X"0F",X"FF",X"FF",X"11",X"F0",X"FF",X"FF",X"F4",X"F0",X"FF",X"FF",
		X"F4",X"F0",X"FF",X"FF",X"11",X"F0",X"FF",X"FF",X"F4",X"F0",X"FF",X"FF",X"F4",X"F0",X"FF",X"FF",
		X"F4",X"F0",X"FF",X"FF",X"11",X"F0",X"FF",X"FF",X"F4",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"FF",X"FF",X"FF",X"78",X"9F",X"FF",X"FF",X"78",X"9F",X"FF",X"FF",X"F9",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AC",X"CC",X"CC",X"CC",X"A2",X"CC",X"CC",X"22",X"A2",X"C2",X"22",X"32",
		X"E2",X"22",X"23",X"32",X"E2",X"22",X"32",X"33",X"E2",X"C2",X"22",X"33",X"E2",X"C2",X"22",X"32",
		X"E2",X"C2",X"2C",X"3C",X"EC",X"CC",X"CC",X"CC",X"88",X"88",X"00",X"00",X"EE",X"E0",X"0E",X"EE",
		X"EE",X"E0",X"00",X"EE",X"EE",X"E0",X"0E",X"00",X"88",X"88",X"88",X"88",X"AA",X"AA",X"A7",X"AA",
		X"AA",X"AA",X"AA",X"97",X"CC",X"AC",X"CA",X"97",X"CC",X"AC",X"CA",X"97",X"33",X"32",X"2A",X"97",
		X"22",X"F2",X"2A",X"97",X"33",X"32",X"CA",X"97",X"22",X"F3",X"2A",X"97",X"22",X"A3",X"2A",X"97",
		X"33",X"32",X"2A",X"97",X"CC",X"AC",X"CA",X"97",X"88",X"80",X"88",X"88",X"0E",X"E0",X"EE",X"E8",
		X"0E",X"E0",X"EE",X"E8",X"0E",X"E0",X"EE",X"E8",X"88",X"88",X"88",X"88",X"77",X"AA",X"AA",X"AA",
		X"F9",X"FF",X"FF",X"9F",X"79",X"FF",X"FF",X"9F",X"79",X"77",X"11",X"9F",X"11",X"77",X"77",X"9F",
		X"11",X"71",X"77",X"1F",X"19",X"11",X"11",X"9F",X"17",X"71",X"77",X"FF",X"19",X"91",X"99",X"9F",
		X"11",X"77",X"33",X"FF",X"11",X"99",X"39",X"9F",X"77",X"77",X"37",X"FF",X"99",X"99",X"99",X"99",
		X"77",X"73",X"33",X"7F",X"93",X"93",X"99",X"99",X"73",X"73",X"77",X"7F",X"77",X"77",X"77",X"7F",
		X"CC",X"CC",X"AA",X"77",X"CC",X"CC",X"AC",X"77",X"44",X"4C",X"A4",X"77",X"44",X"4C",X"A4",X"77",
		X"44",X"4C",X"A4",X"77",X"44",X"4C",X"A4",X"77",X"44",X"4C",X"A4",X"77",X"44",X"4C",X"AA",X"77",
		X"4C",X"CC",X"A4",X"77",X"CC",X"CC",X"A4",X"99",X"99",X"99",X"A4",X"88",X"77",X"77",X"A4",X"88",
		X"77",X"77",X"AC",X"88",X"77",X"77",X"AD",X"88",X"88",X"88",X"CC",X"CC",X"66",X"66",X"66",X"66",
		X"88",X"88",X"88",X"FF",X"77",X"77",X"BB",X"FF",X"82",X"77",X"BE",X"FF",X"72",X"77",X"BB",X"FF",
		X"72",X"77",X"FF",X"CF",X"F3",X"77",X"F8",X"7C",X"33",X"77",X"B8",X"77",X"33",X"B7",X"B8",X"99",
		X"E3",X"BF",X"BB",X"FF",X"33",X"BB",X"BB",X"77",X"33",X"EB",X"BB",X"77",X"33",X"BB",X"BE",X"77",
		X"33",X"BB",X"BB",X"77",X"33",X"FB",X"BB",X"77",X"33",X"77",X"B7",X"77",X"E3",X"77",X"A7",X"77",
		X"80",X"80",X"88",X"88",X"55",X"5F",X"44",X"C3",X"5D",X"57",X"4D",X"A3",X"55",X"57",X"44",X"77",
		X"55",X"F4",X"F4",X"77",X"55",X"44",X"2F",X"77",X"55",X"44",X"2C",X"46",X"5D",X"44",X"22",X"44",
		X"55",X"4D",X"22",X"D4",X"55",X"24",X"22",X"44",X"55",X"22",X"A2",X"44",X"55",X"22",X"4F",X"44",
		X"55",X"22",X"44",X"47",X"55",X"22",X"44",X"77",X"55",X"22",X"44",X"77",X"5D",X"22",X"24",X"77",
		X"FC",X"CF",X"FA",X"CC",X"FC",X"CF",X"F7",X"CC",X"FC",X"CF",X"F7",X"CC",X"FC",X"CF",X"F7",X"CC",
		X"FC",X"CF",X"F7",X"22",X"FC",X"CF",X"F7",X"22",X"FC",X"2F",X"F7",X"22",X"FC",X"2F",X"F7",X"22",
		X"FC",X"2F",X"F7",X"22",X"F2",X"2F",X"FF",X"22",X"F2",X"2F",X"F7",X"22",X"F2",X"2F",X"F7",X"22",
		X"F2",X"2F",X"F7",X"22",X"F2",X"2F",X"F7",X"77",X"F2",X"2F",X"FA",X"22",X"F2",X"2F",X"F7",X"77",
		X"CA",X"AA",X"CC",X"A7",X"CA",X"CC",X"CC",X"A7",X"2A",X"22",X"22",X"A7",X"2A",X"22",X"22",X"A7",
		X"2A",X"22",X"22",X"A7",X"2A",X"22",X"22",X"A7",X"2A",X"22",X"22",X"A7",X"2A",X"AA",X"2C",X"A7",
		X"CA",X"22",X"CC",X"A7",X"CA",X"22",X"CC",X"99",X"9A",X"22",X"99",X"88",X"77",X"22",X"77",X"88",
		X"77",X"CC",X"77",X"88",X"77",X"AA",X"77",X"88",X"88",X"CC",X"88",X"CC",X"66",X"66",X"66",X"66",
		X"F2",X"2F",X"F7",X"22",X"F2",X"2F",X"F7",X"22",X"F2",X"2F",X"F7",X"22",X"F2",X"2F",X"F7",X"22",
		X"F2",X"2F",X"F7",X"22",X"F2",X"2F",X"F7",X"77",X"F2",X"2F",X"F7",X"22",X"FF",X"F2",X"F7",X"22",
		X"FF",X"FF",X"F7",X"22",X"F2",X"2F",X"FF",X"22",X"FA",X"ED",X"F7",X"22",X"F7",X"89",X"F7",X"22",
		X"F7",X"89",X"F7",X"77",X"F7",X"89",X"F7",X"CC",X"7C",X"89",X"77",X"CC",X"66",X"66",X"66",X"66",
		X"7F",X"12",X"22",X"19",X"71",X"22",X"22",X"1F",X"1F",X"11",X"11",X"17",X"7F",X"C2",X"22",X"77",
		X"94",X"CC",X"C2",X"97",X"FF",X"EE",X"EE",X"F7",X"99",X"44",X"44",X"47",X"77",X"77",X"77",X"44",
		X"FF",X"22",X"44",X"47",X"7F",X"24",X"22",X"47",X"7F",X"42",X"22",X"47",X"74",X"22",X"22",X"47",
		X"4F",X"44",X"44",X"49",X"7F",X"22",X"2E",X"FF",X"7F",X"22",X"22",X"F7",X"7F",X"22",X"22",X"F7",
		X"7E",X"77",X"E7",X"99",X"7E",X"77",X"E7",X"FF",X"11",X"77",X"E7",X"7F",X"7E",X"77",X"E7",X"7F",
		X"7E",X"77",X"E7",X"7F",X"7E",X"77",X"E7",X"7F",X"99",X"99",X"99",X"7F",X"74",X"77",X"77",X"7F",
		X"74",X"77",X"E7",X"7F",X"7E",X"77",X"E7",X"7F",X"7E",X"77",X"E7",X"7F",X"7E",X"77",X"E7",X"7F",
		X"44",X"77",X"E7",X"9F",X"7E",X"77",X"E7",X"FF",X"7E",X"77",X"E7",X"77",X"7E",X"77",X"E7",X"77",
		X"7E",X"77",X"E7",X"99",X"7E",X"77",X"E7",X"FF",X"7E",X"77",X"E7",X"7F",X"70",X"77",X"E7",X"7F",
		X"70",X"77",X"E7",X"7F",X"7E",X"77",X"E7",X"7F",X"99",X"99",X"99",X"7F",X"77",X"77",X"77",X"7F",
		X"00",X"77",X"E7",X"7F",X"7E",X"77",X"E7",X"7F",X"7E",X"77",X"E7",X"7F",X"7E",X"77",X"E7",X"7F",
		X"7A",X"77",X"E7",X"9F",X"71",X"77",X"E7",X"FF",X"71",X"77",X"E7",X"77",X"7E",X"77",X"E7",X"77",
		X"70",X"22",X"22",X"79",X"7F",X"22",X"22",X"77",X"7F",X"00",X"00",X"07",X"7F",X"22",X"22",X"00",
		X"9F",X"CC",X"00",X"07",X"FF",X"E0",X"EE",X"07",X"99",X"07",X"79",X"07",X"70",X"77",X"77",X"07",
		X"0F",X"00",X"00",X"07",X"7F",X"22",X"22",X"77",X"71",X"22",X"22",X"77",X"7F",X"22",X"22",X"77",
		X"7F",X"11",X"11",X"19",X"7F",X"22",X"2A",X"11",X"7F",X"22",X"11",X"17",X"7F",X"21",X"22",X"17",
		X"A8",X"F7",X"8F",X"FF",X"88",X"F7",X"8F",X"FF",X"88",X"66",X"66",X"66",X"88",X"77",X"77",X"76",
		X"88",X"37",X"37",X"76",X"8F",X"37",X"37",X"76",X"88",X"77",X"37",X"76",X"88",X"37",X"73",X"36",
		X"88",X"77",X"77",X"73",X"8F",X"33",X"33",X"36",X"99",X"F8",X"8F",X"FF",X"9F",X"F8",X"8F",X"FF",
		X"F9",X"FE",X"8F",X"FF",X"99",X"ED",X"8F",X"FF",X"99",X"DD",X"AF",X"FF",X"99",X"DD",X"AF",X"FF",
		X"77",X"33",X"77",X"77",X"77",X"93",X"77",X"77",X"47",X"33",X"77",X"77",X"47",X"9F",X"77",X"77",
		X"47",X"33",X"77",X"77",X"74",X"93",X"77",X"77",X"74",X"33",X"77",X"77",X"77",X"9F",X"77",X"77",
		X"74",X"33",X"77",X"77",X"74",X"93",X"77",X"77",X"74",X"33",X"77",X"77",X"74",X"9F",X"77",X"77",
		X"74",X"33",X"77",X"77",X"44",X"9F",X"77",X"77",X"44",X"00",X"FF",X"FF",X"77",X"9F",X"77",X"77",
		X"FF",X"FF",X"FF",X"BB",X"CC",X"FF",X"11",X"FF",X"77",X"CC",X"FF",X"11",X"77",X"77",X"FF",X"FF",
		X"77",X"99",X"97",X"FF",X"77",X"88",X"87",X"11",X"77",X"88",X"11",X"FF",X"77",X"8F",X"19",X"99",
		X"99",X"8F",X"F1",X"8F",X"88",X"8F",X"F8",X"8F",X"88",X"8F",X"F8",X"11",X"FF",X"FF",X"FF",X"FF",
		X"8B",X"B8",X"8B",X"B8",X"9B",X"B9",X"9B",X"B9",X"8B",X"B8",X"8B",X"B8",X"FF",X"FF",X"FF",X"FF",
		X"11",X"1C",X"11",X"88",X"11",X"11",X"11",X"88",X"C1",X"11",X"11",X"8F",X"11",X"11",X"11",X"88",
		X"11",X"11",X"11",X"88",X"CC",X"CC",X"CC",X"88",X"99",X"99",X"99",X"88",X"F8",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"F8",X"88",X"88",X"88",X"C8",X"88",X"FF",X"6F",X"FF",X"FF",
		X"66",X"66",X"66",X"66",X"66",X"88",X"66",X"66",X"66",X"76",X"66",X"66",X"66",X"66",X"66",X"66",
		X"FF",X"FF",X"FF",X"FF",X"77",X"77",X"77",X"77",X"CC",X"CC",X"CC",X"77",X"CC",X"CC",X"CC",X"77",
		X"CC",X"CC",X"CC",X"77",X"CC",X"CC",X"CC",X"77",X"11",X"11",X"CC",X"77",X"11",X"11",X"CC",X"77",
		X"11",X"11",X"11",X"88",X"11",X"11",X"11",X"88",X"11",X"11",X"11",X"88",X"11",X"C1",X"11",X"88",
		X"C1",X"1C",X"11",X"88",X"1C",X"11",X"11",X"88",X"11",X"11",X"C1",X"88",X"11",X"11",X"1C",X"88",
		X"FF",X"FF",X"FF",X"FF",X"BB",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"FF",X"1F",X"FB",X"FF",X"FF",
		X"F1",X"99",X"BB",X"FF",X"F8",X"18",X"77",X"FF",X"98",X"18",X"11",X"FF",X"88",X"18",X"17",X"1F",
		X"88",X"18",X"17",X"FF",X"81",X"18",X"17",X"1F",X"18",X"88",X"11",X"1F",X"FF",X"FF",X"FF",X"FF",
		X"B8",X"8B",X"B8",X"87",X"B9",X"9B",X"B9",X"97",X"B8",X"8B",X"B8",X"87",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"33",X"FF",X"FF",X"FF",X"3F",X"FF",X"FF",X"FF",X"3F",X"FF",
		X"FF",X"3F",X"3F",X"FF",X"33",X"FF",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"11",X"1F",X"FF",X"FF",
		X"AA",X"FF",X"FF",X"FF",X"11",X"FF",X"FF",X"FF",X"E1",X"1F",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",
		X"77",X"AA",X"6F",X"DD",X"C7",X"AF",X"7F",X"ED",X"C7",X"FF",X"7C",X"6E",X"C7",X"F6",X"7F",X"7E",
		X"27",X"FF",X"7C",X"7F",X"27",X"FF",X"7F",X"7F",X"27",X"FF",X"7C",X"CF",X"27",X"FF",X"7F",X"7F",
		X"77",X"AE",X"7C",X"7E",X"77",X"AF",X"7A",X"7A",X"77",X"FF",X"7F",X"AA",X"7C",X"FF",X"AA",X"AA",
		X"CF",X"F6",X"AA",X"AA",X"FF",X"66",X"AA",X"2A",X"FF",X"6C",X"EE",X"EA",X"FF",X"66",X"66",X"66",
		X"9E",X"7C",X"79",X"88",X"9E",X"7C",X"79",X"88",X"9E",X"7C",X"79",X"8F",X"9E",X"72",X"79",X"8C",
		X"9E",X"72",X"79",X"F8",X"9E",X"77",X"79",X"C8",X"9E",X"77",X"79",X"87",X"9E",X"77",X"79",X"C7",
		X"9E",X"66",X"69",X"FF",X"9E",X"66",X"69",X"CF",X"9E",X"66",X"69",X"7C",X"9E",X"66",X"69",X"FF",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"76",X"66",X"A6",X"66",X"66",X"66",X"66",X"66",X"67",
		X"77",X"8F",X"88",X"88",X"77",X"8F",X"99",X"88",X"7A",X"FC",X"F9",X"88",X"7A",X"7C",X"F9",X"F8",
		X"7A",X"7C",X"79",X"88",X"7A",X"7C",X"79",X"88",X"7A",X"7C",X"79",X"88",X"9A",X"7C",X"79",X"88",
		X"9A",X"7C",X"79",X"88",X"9A",X"7C",X"79",X"8F",X"9A",X"EE",X"79",X"88",X"FA",X"7C",X"79",X"F8",
		X"CA",X"7C",X"79",X"88",X"9A",X"7C",X"79",X"F8",X"9A",X"7C",X"79",X"88",X"9A",X"7C",X"79",X"88",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"CC",X"CC",X"CC",X"C9",X"CC",X"CC",X"CC",X"99",
		X"77",X"77",X"77",X"99",X"EE",X"EE",X"EE",X"9D",X"EE",X"EE",X"EE",X"D9",X"EE",X"EE",X"EE",X"9D",
		X"EE",X"EE",X"EE",X"D9",X"EE",X"EE",X"EE",X"9D",X"EE",X"EE",X"EE",X"D9",X"EE",X"EE",X"EE",X"99",
		X"EE",X"EE",X"EE",X"99",X"EE",X"EE",X"EE",X"99",X"77",X"77",X"77",X"9F",X"FF",X"FF",X"FF",X"FF",
		X"77",X"7F",X"7F",X"F7",X"77",X"7F",X"7F",X"F7",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"77",X"77",X"77",X"77",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"77",X"77",X"77",X"77",X"FF",X"FF",X"FF",X"FF",
		X"9F",X"6E",X"FF",X"FF",X"9F",X"6E",X"FF",X"FF",X"F6",X"6F",X"FF",X"FF",X"F6",X"EF",X"FF",X"FF",
		X"F6",X"EF",X"FF",X"FF",X"66",X"FF",X"FF",X"FF",X"66",X"FF",X"FF",X"FF",X"67",X"FF",X"FF",X"FF",
		X"66",X"FF",X"FF",X"FF",X"66",X"FF",X"FF",X"FF",X"66",X"FF",X"FF",X"FF",X"66",X"FF",X"FF",X"FF",
		X"66",X"FF",X"FF",X"FF",X"66",X"FF",X"FF",X"FF",X"66",X"FF",X"FF",X"FF",X"66",X"FF",X"FF",X"FF",
		X"99",X"F6",X"6F",X"FF",X"99",X"F6",X"DF",X"FF",X"99",X"F6",X"DF",X"FF",X"99",X"66",X"FF",X"FF",
		X"99",X"66",X"FF",X"FF",X"99",X"66",X"FF",X"FF",X"99",X"66",X"FF",X"FF",X"99",X"66",X"FF",X"FF",
		X"99",X"66",X"FF",X"FF",X"99",X"66",X"FF",X"FF",X"99",X"66",X"FF",X"FF",X"99",X"66",X"FF",X"FF",
		X"99",X"66",X"FF",X"FF",X"99",X"66",X"FF",X"FF",X"99",X"66",X"FF",X"FF",X"9F",X"66",X"FF",X"FF",
		X"44",X"44",X"44",X"88",X"44",X"44",X"44",X"88",X"C4",X"44",X"44",X"88",X"4C",X"44",X"44",X"88",
		X"44",X"44",X"44",X"88",X"CC",X"CC",X"CC",X"88",X"99",X"99",X"99",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",X"FF",X"FF",X"FF",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"FF",X"FF",X"FF",X"FF",X"77",X"77",X"77",X"77",X"CC",X"CC",X"CC",X"77",X"CC",X"CC",X"CC",X"77",
		X"CC",X"CC",X"CC",X"77",X"CC",X"CC",X"CC",X"77",X"44",X"44",X"CC",X"77",X"44",X"44",X"CC",X"77",
		X"44",X"44",X"44",X"88",X"44",X"44",X"44",X"88",X"C4",X"4C",X"44",X"88",X"4C",X"44",X"44",X"88",
		X"C4",X"44",X"C4",X"88",X"4C",X"44",X"4C",X"88",X"44",X"44",X"44",X"88",X"44",X"44",X"44",X"88",
		X"7E",X"77",X"E7",X"99",X"7E",X"77",X"E7",X"FF",X"7E",X"77",X"E7",X"7F",X"7E",X"77",X"E7",X"7F",
		X"7E",X"77",X"E7",X"7F",X"7E",X"77",X"E7",X"7F",X"99",X"99",X"99",X"7F",X"77",X"77",X"77",X"7F",
		X"7E",X"77",X"E7",X"7F",X"7E",X"77",X"E7",X"7F",X"7E",X"77",X"E7",X"7F",X"7E",X"77",X"E7",X"7F",
		X"7E",X"77",X"E7",X"9F",X"7E",X"77",X"E7",X"FF",X"7E",X"77",X"E7",X"77",X"7E",X"77",X"E7",X"77",
		X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FD",X"FF",X"DF",
		X"78",X"FF",X"DD",X"FD",X"78",X"FD",X"DA",X"FF",X"AA",X"FF",X"DA",X"FF",X"77",X"FF",X"DA",X"DA",
		X"77",X"FF",X"FA",X"DA",X"78",X"FF",X"FA",X"FA",X"78",X"FF",X"FA",X"FA",X"78",X"FF",X"FA",X"FA",
		X"78",X"FF",X"FA",X"FA",X"78",X"AF",X"FA",X"FA",X"78",X"FF",X"FA",X"FF",X"78",X"FF",X"FF",X"FF",
		X"22",X"CA",X"CC",X"CC",X"88",X"FA",X"29",X"22",X"88",X"FA",X"29",X"22",X"88",X"FA",X"29",X"22",
		X"88",X"FA",X"29",X"C2",X"88",X"FA",X"29",X"C2",X"88",X"FA",X"C9",X"C2",X"AA",X"CA",X"CA",X"AA",
		X"99",X"FA",X"26",X"66",X"88",X"FA",X"28",X"79",X"88",X"FA",X"C8",X"79",X"88",X"FA",X"C8",X"79",
		X"88",X"FA",X"E8",X"79",X"88",X"FA",X"E8",X"79",X"77",X"CC",X"C7",X"77",X"66",X"66",X"66",X"66",
		X"EE",X"AA",X"AA",X"89",X"AA",X"AA",X"AF",X"89",X"EE",X"AF",X"AF",X"F9",X"CF",X"FF",X"EF",X"F7",
		X"FC",X"FF",X"EF",X"9F",X"CF",X"CF",X"FF",X"6F",X"FC",X"CF",X"FF",X"87",X"CF",X"CF",X"FF",X"89",
		X"AA",X"AE",X"AA",X"89",X"AA",X"AA",X"AA",X"88",X"AA",X"AA",X"EE",X"98",X"AA",X"AA",X"CC",X"CC",
		X"AA",X"A2",X"CC",X"CC",X"A2",X"AA",X"CC",X"CC",X"2E",X"EE",X"CC",X"66",X"66",X"66",X"66",X"66",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"FF",X"FF",X"FF",
		X"AA",X"EF",X"FF",X"FF",X"FF",X"ED",X"FF",X"FF",X"EE",X"ED",X"FF",X"FF",X"EE",X"ED",X"EE",X"F8",
		X"EE",X"ED",X"AA",X"86",X"FF",X"ED",X"EA",X"F7",X"EE",X"ED",X"EA",X"F8",X"EE",X"ED",X"AA",X"98",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"FF",X"FF",X"FF",X"FE",X"DF",
		X"FA",X"FF",X"FE",X"DD",X"88",X"DF",X"FE",X"DD",X"88",X"DD",X"EE",X"DD",X"FF",X"DD",X"FE",X"DD",
		X"AC",X"CC",X"AC",X"CC",X"AC",X"CC",X"AC",X"CC",X"A2",X"C2",X"A2",X"C2",X"A2",X"C2",X"A2",X"22",
		X"A2",X"C2",X"A2",X"22",X"A2",X"22",X"A2",X"22",X"A2",X"22",X"A2",X"AA",X"A2",X"CC",X"A2",X"22",
		X"A2",X"CC",X"A2",X"22",X"A2",X"22",X"A2",X"22",X"99",X"99",X"99",X"22",X"77",X"77",X"77",X"CC",
		X"99",X"99",X"97",X"CC",X"77",X"77",X"97",X"AA",X"77",X"77",X"97",X"CC",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"66",X"66",X"CC",X"76",X"66",X"6C",X"CC",X"66",X"66",X"CC",X"CC",X"66",
		X"66",X"EE",X"EE",X"66",X"EE",X"EF",X"FF",X"EE",X"EE",X"FF",X"FF",X"EE",X"9F",X"EE",X"EE",X"FF",
		X"FF",X"FF",X"FF",X"69",X"FF",X"FF",X"FF",X"99",X"FF",X"F5",X"FF",X"FF",X"FF",X"DD",X"FF",X"FF",
		X"FF",X"DD",X"FF",X"FF",X"FD",X"53",X"FF",X"FF",X"5D",X"DA",X"FF",X"FF",X"FD",X"AB",X"FF",X"FF",
		X"66",X"66",X"66",X"66",X"66",X"66",X"CC",X"76",X"66",X"6C",X"CC",X"66",X"66",X"CC",X"CC",X"66",
		X"66",X"EE",X"EE",X"66",X"E5",X"EF",X"FF",X"EE",X"5E",X"FF",X"FF",X"EE",X"EE",X"5E",X"EE",X"FF",
		X"E5",X"3F",X"FF",X"69",X"E5",X"33",X"FF",X"99",X"EE",X"5F",X"FF",X"FF",X"5E",X"ED",X"FF",X"FF",
		X"F5",X"EE",X"FF",X"FF",X"FE",X"AA",X"FF",X"FF",X"FA",X"AB",X"FF",X"FF",X"FF",X"AA",X"FF",X"FF",
		X"66",X"D5",X"66",X"66",X"63",X"DD",X"CC",X"76",X"33",X"5D",X"CC",X"66",X"65",X"DD",X"CC",X"66",
		X"B6",X"D5",X"EE",X"66",X"EE",X"FF",X"BF",X"EE",X"BE",X"FF",X"FF",X"EE",X"FB",X"9E",X"EE",X"FF",
		X"89",X"79",X"FF",X"69",X"F9",X"17",X"FF",X"99",X"FF",X"77",X"FF",X"FF",X"FF",X"F6",X"FF",X"FF",
		X"FF",X"F6",X"FF",X"FF",X"FA",X"F6",X"FF",X"FF",X"FA",X"67",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"CC",X"CC",X"CC",X"CC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"CC",X"CC",X"CC",X"CC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"FF",X"FE",X"FE",X"FF",X"FF",X"ED",X"DD",X"DE",X"FE",X"DD",
		X"EE",X"ED",X"ED",X"DD",X"DD",X"7D",X"DD",X"DD",X"DD",X"7D",X"DD",X"DD",X"DD",X"7D",X"DD",X"DD",
		X"FA",X"DD",X"AF",X"F7",X"FA",X"DA",X"AF",X"F7",X"FA",X"DA",X"AF",X"F7",X"FA",X"DA",X"FF",X"A7",
		X"FA",X"AA",X"FF",X"A7",X"FF",X"FF",X"FF",X"A7",X"FF",X"FF",X"FF",X"A7",X"FF",X"FF",X"FF",X"A7",
		X"FF",X"FF",X"FF",X"A7",X"FF",X"FF",X"FF",X"A7",X"FF",X"FF",X"FF",X"A7",X"FF",X"FF",X"FF",X"A7",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"DD",X"C7",X"CC",X"7C",X"DD",X"C7",X"CC",X"7C",X"DD",X"C7",X"CC",X"7C",X"FF",X"77",X"CC",X"7C",
		X"F7",X"77",X"CC",X"7C",X"F7",X"7C",X"CC",X"7C",X"F7",X"7C",X"CC",X"7C",X"F7",X"CC",X"CC",X"7C",
		X"F7",X"CC",X"CC",X"7C",X"F7",X"CC",X"CC",X"7C",X"F7",X"CC",X"CC",X"7C",X"F7",X"CC",X"CC",X"7C",
		X"F7",X"CC",X"CC",X"7C",X"F7",X"CC",X"CC",X"7C",X"F7",X"CC",X"CC",X"7C",X"F7",X"CC",X"CC",X"7C",
		X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"EE",X"FF",X"FF",X"EF",X"EE",X"FF",X"FF",X"FE",X"EA",
		X"FF",X"EF",X"DD",X"AA",X"FF",X"FF",X"DF",X"FF",X"FE",X"FE",X"DE",X"FF",X"EE",X"ED",X"DD",X"FF",
		X"EE",X"DD",X"AA",X"FF",X"EE",X"DD",X"FF",X"FF",X"DD",X"DD",X"AF",X"FF",X"DD",X"DD",X"AF",X"FF",
		X"DD",X"DD",X"AF",X"FF",X"AA",X"DD",X"AF",X"FF",X"FF",X"DD",X"AF",X"FF",X"FF",X"DD",X"AF",X"FF",
		X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"C7",X"FF",X"FF",X"FF",X"C7",
		X"FF",X"FF",X"FF",X"C7",X"FF",X"FF",X"FF",X"C7",X"FF",X"FF",X"F8",X"C7",X"FF",X"FF",X"87",X"C7",
		X"FF",X"FF",X"7C",X"C7",X"FF",X"FF",X"CC",X"C7",X"FF",X"FF",X"CC",X"C7",X"FF",X"FE",X"CC",X"C7",
		X"FF",X"E7",X"CC",X"C7",X"FE",X"F7",X"CC",X"C7",X"EE",X"E7",X"CC",X"C7",X"DD",X"77",X"CC",X"C7",
		X"C7",X"77",X"CC",X"C7",X"C7",X"77",X"CC",X"C7",X"77",X"77",X"CC",X"C7",X"77",X"77",X"C7",X"C7",
		X"77",X"77",X"C7",X"C7",X"77",X"77",X"67",X"C7",X"77",X"77",X"77",X"C7",X"77",X"77",X"77",X"77",
		X"77",X"88",X"77",X"77",X"77",X"87",X"77",X"77",X"7F",X"87",X"77",X"77",X"7F",X"87",X"77",X"77",
		X"AF",X"87",X"77",X"77",X"AA",X"AA",X"77",X"77",X"AA",X"AA",X"AA",X"77",X"AA",X"AA",X"AA",X"AA",
		X"11",X"11",X"11",X"99",X"FF",X"FF",X"FF",X"99",X"FB",X"BB",X"FF",X"99",X"FF",X"BF",X"FF",X"99",
		X"FF",X"FF",X"FF",X"99",X"FF",X"BB",X"FF",X"99",X"FF",X"FF",X"FF",X"99",X"11",X"11",X"11",X"99",
		X"FF",X"FF",X"88",X"99",X"F1",X"FF",X"88",X"99",X"1F",X"F8",X"88",X"99",X"FF",X"88",X"88",X"99",
		X"FF",X"88",X"88",X"99",X"FF",X"88",X"87",X"99",X"11",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"F1",X"11",X"11",X"11",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"BF",X"FF",X"FB",X"BB",X"FB",
		X"FF",X"FB",X"BF",X"BF",X"FF",X"FF",X"BF",X"FF",X"1F",X"FF",X"FF",X"FF",X"71",X"11",X"F1",X"F1",
		X"77",X"FF",X"FF",X"F1",X"77",X"88",X"FF",X"F1",X"78",X"88",X"FF",X"F1",X"88",X"88",X"FF",X"F1",
		X"88",X"88",X"FF",X"F1",X"88",X"88",X"FF",X"F1",X"99",X"99",X"11",X"F1",X"99",X"99",X"88",X"88",
		X"22",X"A2",X"27",X"67",X"22",X"A2",X"27",X"F7",X"22",X"A2",X"27",X"77",X"22",X"A2",X"27",X"77",
		X"22",X"A2",X"27",X"77",X"22",X"A2",X"27",X"77",X"22",X"A2",X"27",X"77",X"CC",X"AC",X"C8",X"67",
		X"88",X"88",X"88",X"67",X"22",X"A2",X"27",X"F7",X"22",X"A2",X"27",X"77",X"22",X"A2",X"27",X"77",
		X"22",X"A2",X"27",X"77",X"22",X"A2",X"27",X"77",X"22",X"A2",X"27",X"77",X"22",X"A2",X"27",X"67",
		X"98",X"99",X"87",X"7F",X"98",X"99",X"87",X"7F",X"98",X"99",X"87",X"7F",X"AA",X"A2",X"AA",X"A2",
		X"EE",X"22",X"2E",X"22",X"EE",X"EE",X"EE",X"EE",X"1E",X"EE",X"EE",X"EE",X"E1",X"1E",X"EE",X"EE",
		X"1E",X"E1",X"EE",X"EE",X"11",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"E3",X"1E",X"EE",X"EE",
		X"E3",X"EE",X"EE",X"EE",X"A3",X"AA",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"77",X"77",X"77",X"77",
		X"FF",X"99",X"FF",X"FF",X"F9",X"55",X"F9",X"FF",X"F5",X"55",X"F5",X"99",X"F5",X"55",X"F5",X"55",
		X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"99",X"F7",X"55",X"F7",X"99",X"F7",X"79",
		X"F7",X"55",X"F7",X"79",X"F5",X"55",X"F5",X"79",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",
		X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"55",X"F5",X"99",X"F7",X"55",X"F7",X"99",X"F7",X"79",
		X"FC",X"F2",X"22",X"AA",X"FC",X"F2",X"22",X"22",X"FC",X"F2",X"2C",X"22",X"FC",X"F2",X"2C",X"2C",
		X"FC",X"F2",X"2C",X"2C",X"FC",X"F2",X"2C",X"2C",X"FC",X"F2",X"2C",X"2C",X"FC",X"F2",X"2C",X"AA",
		X"FC",X"F2",X"2C",X"2C",X"FC",X"FC",X"CC",X"CC",X"FC",X"F2",X"22",X"22",X"FC",X"F2",X"22",X"22",
		X"F2",X"F2",X"22",X"22",X"CC",X"CC",X"CC",X"AA",X"77",X"77",X"77",X"CC",X"66",X"66",X"66",X"66",
		X"67",X"FF",X"F7",X"F2",X"27",X"FF",X"F7",X"F2",X"77",X"FE",X"F7",X"F2",X"77",X"FE",X"F7",X"F2",
		X"77",X"FE",X"F7",X"F2",X"77",X"FE",X"F7",X"F2",X"77",X"FF",X"F7",X"F2",X"77",X"FF",X"F7",X"F2",
		X"77",X"FF",X"F7",X"F2",X"77",X"FF",X"F7",X"F7",X"77",X"FF",X"F7",X"F7",X"76",X"FF",X"CF",X"FC",
		X"6F",X"F6",X"FC",X"FF",X"FF",X"66",X"CC",X"FC",X"FF",X"66",X"66",X"66",X"FF",X"66",X"66",X"66",
		X"77",X"67",X"77",X"77",X"77",X"F6",X"99",X"F9",X"77",X"F8",X"88",X"88",X"77",X"FF",X"FC",X"FC",
		X"77",X"FF",X"F2",X"F2",X"77",X"FF",X"F2",X"F2",X"77",X"FF",X"F2",X"F2",X"77",X"88",X"8F",X"88",
		X"77",X"99",X"99",X"F9",X"77",X"88",X"88",X"88",X"77",X"EE",X"F7",X"FC",X"77",X"DE",X"F7",X"FC",
		X"77",X"DD",X"F7",X"F2",X"77",X"AA",X"F7",X"F2",X"77",X"FF",X"F7",X"F2",X"77",X"FF",X"F7",X"F2",
		X"77",X"77",X"77",X"77",X"99",X"99",X"99",X"99",X"78",X"88",X"88",X"77",X"99",X"99",X"99",X"99",
		X"78",X"88",X"88",X"77",X"99",X"99",X"99",X"99",X"78",X"88",X"88",X"88",X"99",X"99",X"FF",X"FF",
		X"99",X"99",X"77",X"77",X"78",X"88",X"77",X"77",X"FF",X"FF",X"77",X"77",X"77",X"77",X"77",X"77",
		X"88",X"88",X"88",X"88",X"99",X"99",X"99",X"99",X"88",X"88",X"88",X"88",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"8F",X"FA",X"7F",X"FF",X"8F",X"AA",X"7F",X"FF",X"8F",X"A8",X"7F",X"FF",X"8F",X"A8",X"7F",X"FF",
		X"8F",X"A8",X"8F",X"FF",X"8F",X"88",X"8F",X"FF",X"8F",X"88",X"8F",X"FF",X"8F",X"F8",X"8F",X"FF",
		X"8F",X"F8",X"8F",X"FF",X"8F",X"F8",X"8F",X"FF",X"8F",X"F8",X"8F",X"FF",X"8A",X"F8",X"8F",X"FF",
		X"8A",X"F8",X"8F",X"FF",X"AA",X"F8",X"8F",X"FF",X"AA",X"F8",X"8F",X"FF",X"A8",X"F8",X"8F",X"FF",
		X"88",X"AA",X"AA",X"DD",X"99",X"CA",X"CA",X"CC",X"99",X"CA",X"CA",X"22",X"69",X"2A",X"2A",X"2C",
		X"69",X"2E",X"2A",X"2C",X"C9",X"2E",X"2A",X"2C",X"C9",X"AD",X"AA",X"2C",X"69",X"2D",X"2A",X"77",
		X"C9",X"2D",X"2A",X"CC",X"99",X"2D",X"2A",X"66",X"99",X"2D",X"2A",X"77",X"79",X"DD",X"AA",X"99",
		X"99",X"CC",X"CC",X"99",X"99",X"CC",X"CC",X"99",X"88",X"CC",X"CC",X"77",X"66",X"66",X"66",X"66",
		X"A8",X"F7",X"CA",X"FF",X"88",X"F7",X"2A",X"FF",X"88",X"F7",X"2A",X"FF",X"88",X"F7",X"2A",X"FF",
		X"88",X"F7",X"2A",X"FF",X"88",X"F7",X"2A",X"FF",X"88",X"F7",X"C9",X"FF",X"88",X"F8",X"C9",X"FF",
		X"88",X"F8",X"C7",X"FF",X"89",X"F9",X"97",X"FF",X"99",X"F9",X"7F",X"FF",X"99",X"F9",X"7F",X"FF",
		X"99",X"DD",X"7F",X"FF",X"99",X"DD",X"7F",X"FF",X"99",X"DD",X"AF",X"FF",X"99",X"DD",X"AF",X"FF",
		X"FE",X"2E",X"22",X"FF",X"EE",X"2E",X"22",X"EE",X"7F",X"7F",X"77",X"77",X"7F",X"2F",X"22",X"88",
		X"7F",X"2F",X"22",X"88",X"7F",X"7F",X"77",X"99",X"8F",X"2F",X"22",X"99",X"8F",X"2F",X"22",X"99",
		X"8F",X"7F",X"77",X"99",X"9F",X"2F",X"22",X"99",X"9F",X"2F",X"2C",X"99",X"9F",X"7F",X"77",X"99",
		X"9F",X"CF",X"CC",X"99",X"9F",X"CF",X"CC",X"99",X"9F",X"7F",X"77",X"99",X"9F",X"CF",X"CC",X"DD",
		X"8F",X"88",X"F8",X"FF",X"A8",X"CA",X"8A",X"CC",X"AF",X"CA",X"FA",X"CC",X"AF",X"CA",X"FA",X"22",
		X"AF",X"2A",X"FA",X"22",X"AF",X"2A",X"FA",X"22",X"AF",X"2A",X"FA",X"22",X"AF",X"2A",X"FA",X"AA",
		X"AF",X"2A",X"FA",X"22",X"AF",X"2A",X"FA",X"22",X"AF",X"2A",X"FA",X"22",X"AF",X"CA",X"FA",X"22",
		X"AF",X"2A",X"FA",X"CC",X"AF",X"FA",X"FA",X"AA",X"AC",X"CC",X"CA",X"CC",X"66",X"66",X"66",X"66",
		X"44",X"00",X"77",X"77",X"44",X"F9",X"77",X"77",X"74",X"00",X"77",X"77",X"44",X"F9",X"77",X"77",
		X"44",X"00",X"77",X"77",X"44",X"F9",X"77",X"77",X"74",X"00",X"77",X"77",X"77",X"F9",X"77",X"77",
		X"74",X"00",X"77",X"77",X"74",X"F0",X"77",X"77",X"44",X"00",X"77",X"77",X"44",X"F9",X"77",X"77",
		X"74",X"09",X"77",X"77",X"77",X"F0",X"77",X"77",X"FF",X"00",X"FF",X"FF",X"77",X"F9",X"77",X"77",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"44",X"4F",X"44",X"FF",X"4F",X"FF",X"F4",
		X"FF",X"44",X"FF",X"F4",X"FF",X"4F",X"FF",X"F4",X"FF",X"4F",X"4F",X"F4",X"FF",X"4F",X"FF",X"FF",
		X"FF",X"FF",X"11",X"1F",X"FF",X"FF",X"1F",X"FF",X"FF",X"FF",X"11",X"FF",X"FF",X"FF",X"1F",X"FF",
		X"88",X"88",X"11",X"18",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",
		X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",
		X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DD",X"DD",X"DD",X"DD",
		X"D5",X"55",X"55",X"55",X"AC",X"CC",X"CC",X"CC",X"A5",X"CC",X"CC",X"CC",X"A5",X"55",X"55",X"55",
		X"A5",X"55",X"55",X"55",X"A5",X"55",X"55",X"55",X"A5",X"55",X"55",X"55",X"A5",X"5C",X"55",X"5C",
		X"A5",X"5C",X"55",X"5C",X"A5",X"5C",X"55",X"5C",X"88",X"88",X"88",X"88",X"AA",X"EE",X"EE",X"EE",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"CC",X"CC",X"CC",X"C9",X"CC",X"CC",X"CC",X"99",
		X"77",X"77",X"77",X"99",X"55",X"55",X"55",X"91",X"55",X"55",X"55",X"19",X"55",X"55",X"55",X"90",
		X"33",X"33",X"33",X"09",X"33",X"33",X"33",X"9B",X"33",X"33",X"33",X"B9",X"44",X"44",X"44",X"99",
		X"44",X"44",X"44",X"99",X"44",X"44",X"44",X"99",X"77",X"77",X"77",X"9F",X"FF",X"FF",X"FF",X"FF",
		X"77",X"7F",X"7F",X"F7",X"77",X"7F",X"7F",X"F7",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"77",X"77",X"77",X"77",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"77",X"77",X"77",X"77",X"FF",X"FF",X"FF",X"FF",
		X"22",X"A2",X"27",X"67",X"22",X"A2",X"27",X"F7",X"20",X"AC",X"44",X"77",X"20",X"A0",X"C7",X"77",
		X"20",X"0C",X"27",X"77",X"C0",X"0C",X"27",X"77",X"C0",X"0C",X"27",X"77",X"CC",X"AC",X"C8",X"67",
		X"88",X"88",X"88",X"67",X"C4",X"44",X"44",X"F7",X"4C",X"C4",X"C7",X"77",X"4C",X"A4",X"C7",X"77",
		X"4C",X"A4",X"44",X"77",X"4C",X"A4",X"C7",X"77",X"C4",X"A4",X"44",X"77",X"2C",X"A2",X"C7",X"67",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"4F",X"44",X"FF",X"FF",X"4F",X"44",X"FF",X"FF",
		X"4F",X"44",X"FF",X"FF",X"4F",X"44",X"FF",X"FF",X"4F",X"44",X"FF",X"FF",X"FF",X"44",X"FF",X"FF",
		X"F1",X"4F",X"FF",X"FF",X"1F",X"FF",X"FF",X"FF",X"F1",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"11",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"89",X"89",X"99",X"FF",X"99",X"99",X"97",X"FF",X"99",X"99",X"77",X"FF",
		X"99",X"99",X"7A",X"FF",X"99",X"F8",X"CA",X"FF",X"99",X"F9",X"CA",X"FF",X"FF",X"F9",X"2A",X"FF",
		X"99",X"F9",X"2A",X"FF",X"99",X"F9",X"2A",X"FF",X"99",X"F9",X"2A",X"FF",X"9F",X"F9",X"CA",X"FF",
		X"9F",X"F8",X"C9",X"FF",X"F9",X"F8",X"C9",X"FF",X"F9",X"F8",X"97",X"FF",X"97",X"F7",X"8F",X"FF",
		X"AC",X"CC",X"A8",X"CC",X"AC",X"CC",X"A8",X"CC",X"A2",X"22",X"A8",X"22",X"A2",X"22",X"A9",X"22",
		X"A2",X"22",X"A9",X"22",X"A2",X"C2",X"A9",X"22",X"A2",X"C2",X"A9",X"AA",X"A2",X"CC",X"A9",X"22",
		X"A2",X"CC",X"A9",X"22",X"A2",X"C2",X"A9",X"22",X"AC",X"C2",X"A9",X"22",X"AC",X"CC",X"A9",X"22",
		X"AC",X"CC",X"A9",X"22",X"99",X"99",X"99",X"AA",X"77",X"77",X"79",X"CC",X"66",X"66",X"66",X"66",
		X"55",X"F7",X"7F",X"77",X"55",X"F7",X"7F",X"77",X"75",X"77",X"7F",X"F7",X"75",X"F5",X"5F",X"5F",
		X"75",X"F5",X"5F",X"F7",X"75",X"F5",X"77",X"F7",X"75",X"55",X"75",X"55",X"75",X"FF",X"FF",X"FF",
		X"55",X"FB",X"F7",X"BF",X"5F",X"FB",X"BF",X"BB",X"77",X"F3",X"3F",X"33",X"77",X"F3",X"F7",X"33",
		X"77",X"F3",X"3F",X"33",X"77",X"F4",X"4F",X"44",X"77",X"F4",X"4F",X"44",X"77",X"F4",X"FF",X"44",
		X"77",X"5F",X"77",X"77",X"77",X"5F",X"77",X"77",X"77",X"5F",X"77",X"77",X"55",X"55",X"77",X"77",
		X"55",X"5F",X"77",X"57",X"7F",X"5F",X"77",X"F5",X"55",X"5F",X"F5",X"F5",X"FF",X"FA",X"5F",X"F5",
		X"BB",X"F7",X"55",X"F5",X"BB",X"F7",X"77",X"57",X"3A",X"F7",X"77",X"57",X"3A",X"33",X"77",X"57",
		X"3F",X"33",X"77",X"77",X"4F",X"FF",X"77",X"77",X"4F",X"F7",X"77",X"77",X"4F",X"F7",X"77",X"77",
		X"FF",X"FF",X"FF",X"FF",X"99",X"99",X"F9",X"99",X"7F",X"FF",X"FA",X"77",X"F9",X"9F",X"99",X"88",
		X"8F",X"99",X"99",X"88",X"8F",X"99",X"77",X"99",X"99",X"99",X"88",X"77",X"99",X"99",X"88",X"88",
		X"99",X"F9",X"99",X"88",X"99",X"F7",X"79",X"99",X"77",X"9D",X"99",X"99",X"88",X"99",X"99",X"FF",
		X"99",X"F9",X"99",X"99",X"99",X"8F",X"99",X"F9",X"77",X"8F",X"77",X"FF",X"77",X"97",X"77",X"9F",
		X"FF",X"66",X"66",X"66",X"FF",X"66",X"66",X"66",X"F6",X"66",X"66",X"66",X"F8",X"88",X"88",X"88",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"66",X"66",X"66",X"FF",X"66",X"66",X"66",X"FF",X"66",X"66",X"66",X"FF",X"88",X"88",X"88",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F7",X"99",X"F7",X"79",X"F7",X"99",X"F7",X"79",X"F7",X"99",X"F7",X"79",X"AA",X"A2",X"AA",X"22",
		X"2E",X"22",X"2E",X"22",X"EE",X"EE",X"EE",X"EE",X"EE",X"11",X"E1",X"11",X"EE",X"1E",X"E1",X"EE",
		X"EE",X"11",X"E1",X"E1",X"EE",X"1E",X"E1",X"11",X"EE",X"1E",X"EE",X"EE",X"EE",X"11",X"3E",X"33",
		X"EE",X"EE",X"3E",X"E3",X"AA",X"AA",X"3A",X"A3",X"FF",X"FF",X"FF",X"FF",X"77",X"77",X"77",X"77",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"88",X"88",X"88",X"88",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F7",X"99",X"F7",X"22",X"F7",X"99",X"F7",X"22",X"F7",X"99",X"F7",X"22",X"F7",X"99",X"F7",X"22",
		X"F7",X"99",X"F7",X"22",X"F7",X"99",X"F7",X"22",X"F7",X"99",X"F7",X"22",X"F7",X"99",X"F7",X"22",
		X"F7",X"99",X"F7",X"22",X"F7",X"99",X"FF",X"FF",X"FA",X"EE",X"F7",X"22",X"F8",X"77",X"F7",X"22",
		X"F8",X"77",X"F7",X"FF",X"F8",X"77",X"F7",X"CC",X"CC",X"CC",X"C7",X"CC",X"66",X"66",X"66",X"66",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",
		X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",
		X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"2F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"99",X"FF",X"FF",X"F7",X"55",X"FF",X"FF",X"F7",X"55",
		X"FF",X"FF",X"F7",X"55",X"FF",X"FF",X"F9",X"99",X"FF",X"FF",X"FF",X"88",X"FF",X"FF",X"FF",X"99",
		X"E7",X"DD",X"EE",X"DD",X"F7",X"7D",X"EA",X"EA",X"77",X"E7",X"EA",X"EA",X"F7",X"FF",X"EA",X"EA",
		X"F7",X"CF",X"FA",X"EA",X"99",X"99",X"FA",X"EA",X"88",X"88",X"FF",X"EA",X"99",X"99",X"FC",X"EA",
		X"88",X"88",X"99",X"9A",X"88",X"88",X"88",X"9F",X"77",X"88",X"88",X"89",X"77",X"88",X"78",X"89",
		X"77",X"88",X"77",X"89",X"77",X"88",X"77",X"89",X"77",X"88",X"77",X"77",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"99",X"FF",X"FF",X"FF",X"99",X"F0",X"00",X"0F",X"99",X"90",X"FF",X"FF",X"99",
		X"09",X"FF",X"0F",X"99",X"07",X"FF",X"FF",X"99",X"79",X"00",X"09",X"99",X"97",X"FF",X"97",X"99",
		X"33",X"3F",X"33",X"9F",X"37",X"37",X"33",X"F7",X"33",X"39",X"39",X"77",X"F9",X"99",X"99",X"77",
		X"FF",X"FF",X"FF",X"88",X"99",X"99",X"99",X"99",X"88",X"88",X"88",X"88",X"FF",X"FF",X"FF",X"FF",
		X"88",X"88",X"88",X"F8",X"88",X"A2",X"CC",X"88",X"8F",X"22",X"CC",X"88",X"7F",X"FF",X"FF",X"77",
		X"7F",X"CC",X"CC",X"77",X"7F",X"CC",X"CC",X"77",X"7F",X"CC",X"22",X"77",X"7F",X"CC",X"22",X"77",
		X"7F",X"CC",X"22",X"77",X"7F",X"CC",X"22",X"77",X"7F",X"C2",X"22",X"77",X"7F",X"C2",X"22",X"77",
		X"7F",X"C2",X"22",X"77",X"7F",X"22",X"22",X"77",X"7F",X"22",X"22",X"77",X"7F",X"22",X"22",X"77",
		X"80",X"80",X"88",X"88",X"F8",X"F8",X"22",X"CA",X"88",X"88",X"2C",X"A7",X"77",X"7A",X"FF",X"77",
		X"77",X"7A",X"AC",X"77",X"77",X"7E",X"AC",X"77",X"77",X"7E",X"AC",X"77",X"77",X"7E",X"A2",X"77",
		X"77",X"7E",X"A2",X"77",X"77",X"7E",X"A2",X"77",X"77",X"7E",X"A2",X"77",X"77",X"7E",X"A2",X"77",
		X"77",X"7E",X"A2",X"77",X"77",X"7E",X"A2",X"77",X"77",X"7A",X"A2",X"77",X"77",X"7A",X"A2",X"77",
		X"88",X"76",X"99",X"AA",X"88",X"76",X"99",X"AA",X"78",X"76",X"99",X"A2",X"78",X"76",X"97",X"AA",
		X"88",X"76",X"96",X"EE",X"88",X"76",X"89",X"EE",X"88",X"76",X"89",X"EE",X"88",X"76",X"89",X"EE",
		X"88",X"7F",X"88",X"AA",X"88",X"7C",X"88",X"EE",X"88",X"7C",X"8F",X"EE",X"78",X"76",X"78",X"EE",
		X"F7",X"76",X"F8",X"EE",X"AF",X"76",X"78",X"AA",X"AA",X"F6",X"77",X"66",X"AA",X"A6",X"77",X"66",
		X"AA",X"AA",X"DF",X"AA",X"77",X"77",X"7F",X"77",X"77",X"77",X"7F",X"78",X"77",X"78",X"7F",X"E8",
		X"77",X"78",X"7F",X"E8",X"77",X"88",X"7F",X"E8",X"77",X"87",X"7F",X"A7",X"77",X"87",X"7F",X"A7",
		X"77",X"77",X"7F",X"A7",X"77",X"77",X"7F",X"A7",X"78",X"87",X"7F",X"A7",X"78",X"87",X"7F",X"A7",
		X"78",X"77",X"7F",X"A7",X"88",X"76",X"7F",X"D7",X"87",X"76",X"77",X"77",X"88",X"76",X"99",X"99",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"F7",X"77",X"FF",X"88",X"F7",X"77",
		X"AA",X"88",X"D7",X"FF",X"88",X"88",X"67",X"88",X"88",X"88",X"97",X"88",X"A8",X"A8",X"DF",X"88",
		X"A8",X"A8",X"AF",X"82",X"A8",X"AF",X"86",X"22",X"A7",X"F8",X"86",X"22",X"A7",X"88",X"86",X"82",
		X"F7",X"78",X"86",X"88",X"8F",X"77",X"86",X"88",X"FF",X"77",X"76",X"88",X"77",X"77",X"77",X"77",
		X"FF",X"FE",X"FF",X"DD",X"F1",X"F1",X"1A",X"1F",X"81",X"1F",X"1F",X"AA",X"F1",X"1F",X"A1",X"FF",
		X"F1",X"F1",X"A1",X"1F",X"11",X"FF",X"F1",X"FF",X"8F",X"88",X"88",X"FF",X"87",X"1F",X"81",X"FF",
		X"F1",X"F1",X"81",X"FF",X"F1",X"FF",X"88",X"FF",X"81",X"F8",X"88",X"FF",X"87",X"F8",X"18",X"AF",
		X"88",X"F8",X"F8",X"AA",X"CA",X"CC",X"CC",X"AA",X"CA",X"CC",X"CC",X"CA",X"C9",X"CC",X"CC",X"CC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"FF",
		X"FF",X"FF",X"CF",X"CC",X"FF",X"FF",X"CF",X"DF",X"FF",X"33",X"CF",X"DF",X"FF",X"77",X"77",X"77",
		X"DA",X"FF",X"FF",X"CC",X"DA",X"AA",X"FF",X"CF",X"DA",X"AF",X"DF",X"CC",X"DA",X"AF",X"DD",X"FF",
		X"FF",X"FF",X"DD",X"DD",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"F6",X"6F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"F8",X"FF",X"FF",X"F7",X"66",X"FF",X"AA",X"7F",X"77",X"AA",X"AA",X"FA",X"77",X"AA",
		X"AA",X"E2",X"77",X"CA",X"CC",X"7F",X"77",X"FC",X"CC",X"FF",X"FF",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"FF",X"AA",X"AA",X"AA",X"FF",X"FF",X"CC",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"CF",X"FF",X"FF",X"FF",X"CF",X"FF",X"FF",X"FF",X"FC",X"87",X"FF",X"CC",X"CC",
		X"F8",X"FF",X"CF",X"CC",X"F6",X"FF",X"CF",X"FC",X"86",X"FF",X"CF",X"FC",X"66",X"FF",X"CF",X"FC",
		X"66",X"FF",X"CC",X"CC",X"F2",X"FF",X"FF",X"CF",X"FF",X"FF",X"FF",X"CF",X"DF",X"FF",X"FF",X"FC",
		X"AA",X"A6",X"AA",X"CC",X"AA",X"AA",X"AA",X"CC",X"AA",X"AD",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"EE",X"AA",X"AA",X"AA",X"CE",X"AA",X"AA",X"AA",X"FE",X"AA",X"AA",X"AA",
		X"AF",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EE",X"AA",X"AA",X"AA",X"ED",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"FC",X"CC",X"F6",X"C6",X"CC",X"CC",X"C6",X"C6",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CA",X"CC",X"2C",X"CC",X"AA",X"CC",X"CC",X"CC",X"AA",
		X"CC",X"CC",X"CC",X"CA",X"CC",X"CC",X"CC",X"AA",X"AA",X"88",X"CC",X"AA",X"AA",X"88",X"CC",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"CA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"DA",X"AA",X"AA",X"AA",X"AA",X"DD",X"AA",X"AA",X"66",X"EC",X"CC",X"CC",X"66",X"EC",X"CC",X"FC",
		X"C9",X"CC",X"2C",X"CC",X"C9",X"2E",X"CC",X"CA",X"F9",X"EF",X"FF",X"AA",X"F7",X"CC",X"CC",X"AA",
		X"CC",X"CC",X"CC",X"AA",X"AA",X"CC",X"CA",X"AA",X"AA",X"CC",X"AA",X"AC",X"AA",X"AA",X"AA",X"AC",
		X"AA",X"DD",X"AA",X"CF",X"CA",X"AA",X"AA",X"CF",X"AA",X"AA",X"AA",X"FF",X"AA",X"AE",X"AA",X"FF",
		X"AA",X"AA",X"AA",X"FF",X"AA",X"FF",X"AA",X"FF",X"CC",X"FC",X"C6",X"FF",X"CF",X"CC",X"CC",X"FF",
		X"77",X"FF",X"11",X"1F",X"07",X"77",X"FF",X"F1",X"07",X"70",X"FF",X"F1",X"07",X"70",X"F1",X"F1",
		X"07",X"70",X"FF",X"F1",X"07",X"70",X"11",X"1F",X"07",X"70",X"FF",X"FF",X"07",X"70",X"4F",X"F4",
		X"07",X"70",X"FF",X"4F",X"07",X"70",X"FF",X"4F",X"07",X"70",X"4F",X"4F",X"07",X"70",X"77",X"84",
		X"07",X"70",X"07",X"78",X"07",X"70",X"07",X"78",X"07",X"70",X"07",X"78",X"F2",X"2F",X"F7",X"22",
		X"FF",X"FF",X"99",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"AA",X"6C",X"77",X"FF",X"88",X"C7",X"77",
		X"AA",X"88",X"FF",X"FF",X"88",X"88",X"CC",X"88",X"88",X"88",X"97",X"88",X"A8",X"A8",X"DF",X"88",
		X"A8",X"A8",X"AF",X"82",X"A8",X"AF",X"86",X"22",X"A7",X"F8",X"86",X"22",X"A7",X"88",X"86",X"82",
		X"F7",X"78",X"86",X"88",X"8F",X"77",X"86",X"88",X"FF",X"77",X"76",X"88",X"77",X"77",X"77",X"77",
		X"FF",X"FF",X"AA",X"AA",X"FF",X"FF",X"AA",X"AA",X"FF",X"FF",X"AA",X"AA",X"FF",X"FF",X"CC",X"CC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"DD",X"7D",X"AA",X"AA",X"DD",X"7A",X"FF",X"FA",X"DA",X"7F",X"FF",X"FA",X"DA",X"7F",X"FF",X"FA",
		X"AF",X"7F",X"FF",X"FA",X"AF",X"7F",X"FF",X"FA",X"FF",X"7F",X"FF",X"FF",X"F2",X"7F",X"FF",X"FF",
		X"FF",X"7F",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FC",X"7A",X"AA",X"AA",
		X"FF",X"7A",X"AA",X"AA",X"FF",X"AA",X"AA",X"AA",X"FF",X"FC",X"AA",X"AA",X"FF",X"FF",X"AA",X"AA",
		X"6E",X"66",X"66",X"66",X"6F",X"66",X"66",X"6E",X"66",X"66",X"F6",X"66",X"88",X"88",X"88",X"88",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"99",X"99",X"FF",X"FF",X"77",X"79",X"FF",X"FF",
		X"88",X"F8",X"FF",X"FF",X"88",X"F8",X"FF",X"FF",X"88",X"F8",X"FF",X"FF",X"88",X"FF",X"FF",X"FF",
		X"7F",X"F8",X"FF",X"FF",X"FF",X"F8",X"FF",X"FF",X"9F",X"F8",X"FF",X"FF",X"7F",X"F8",X"FF",X"FF",
		X"79",X"DD",X"AF",X"FF",X"79",X"DD",X"AF",X"FF",X"79",X"DD",X"AF",X"FF",X"79",X"DD",X"AF",X"FF",
		X"79",X"DD",X"AF",X"FF",X"79",X"DD",X"A6",X"FF",X"79",X"DD",X"A6",X"FF",X"66",X"DD",X"A6",X"FF",
		X"AA",X"DD",X"A6",X"FF",X"EE",X"DD",X"A6",X"FF",X"79",X"DD",X"A6",X"FF",X"79",X"DD",X"A6",X"FF",
		X"79",X"DD",X"66",X"FF",X"79",X"DD",X"66",X"FF",X"79",X"DD",X"6D",X"FF",X"99",X"FF",X"6D",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"FF",X"FF",X"99",X"ED",X"FF",X"FF",X"99",X"DD",X"AF",X"FF",X"99",X"DD",X"AF",X"FF",
		X"FF",X"7F",X"77",X"FF",X"FF",X"77",X"77",X"FF",X"FF",X"77",X"A7",X"99",X"F9",X"7F",X"A7",X"99",
		X"89",X"EE",X"A7",X"99",X"89",X"7F",X"A7",X"99",X"89",X"7F",X"A7",X"78",X"89",X"7F",X"A9",X"88",
		X"89",X"7F",X"A9",X"88",X"88",X"7F",X"A9",X"88",X"88",X"7F",X"A9",X"88",X"88",X"FF",X"A9",X"88",
		X"88",X"FF",X"A9",X"88",X"88",X"DE",X"A9",X"88",X"88",X"EE",X"A9",X"88",X"8F",X"99",X"98",X"7F",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"88",X"88",X"88",X"88",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"99",X"99",X"99",X"FF",X"77",X"77",X"77",
		X"99",X"88",X"A6",X"88",X"77",X"88",X"C6",X"88",X"88",X"88",X"AC",X"88",X"8F",X"88",X"AC",X"88",
		X"88",X"88",X"88",X"C8",X"88",X"88",X"88",X"C8",X"99",X"88",X"99",X"88",X"77",X"99",X"77",X"99",
		X"66",X"66",X"66",X"66",X"66",X"66",X"CC",X"76",X"66",X"6C",X"CC",X"66",X"66",X"CC",X"CC",X"66",
		X"66",X"EE",X"EE",X"66",X"EE",X"EF",X"FF",X"EE",X"EE",X"FF",X"FF",X"EE",X"9F",X"EE",X"EE",X"FF",
		X"FF",X"FF",X"FF",X"69",X"FF",X"FF",X"FF",X"99",X"FF",X"FF",X"FF",X"FF",X"FF",X"D5",X"FF",X"FF",
		X"FF",X"DD",X"FF",X"FF",X"FD",X"5D",X"FF",X"FF",X"F5",X"DD",X"FF",X"FF",X"FF",X"D5",X"FF",X"FF",
		X"8C",X"FF",X"FF",X"FF",X"78",X"FF",X"FF",X"FF",X"EF",X"FF",X"FF",X"FF",X"EF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"88",X"88",X"88",X"88",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"99",X"99",X"99",X"99",X"77",X"77",X"77",X"77",
		X"88",X"88",X"88",X"88",X"88",X"AA",X"FF",X"88",X"88",X"AA",X"88",X"88",X"8F",X"CC",X"88",X"88",
		X"FF",X"CC",X"87",X"88",X"88",X"88",X"77",X"98",X"99",X"88",X"99",X"78",X"79",X"99",X"77",X"77",
		X"8F",X"F8",X"FF",X"FF",X"8F",X"F8",X"FF",X"FF",X"8F",X"F8",X"FF",X"FF",X"8F",X"F8",X"FF",X"FF",
		X"8F",X"F8",X"FF",X"FF",X"8F",X"F8",X"FF",X"FF",X"8F",X"F8",X"FF",X"FF",X"8F",X"F8",X"FF",X"FF",
		X"8F",X"F8",X"FF",X"FF",X"8F",X"F8",X"FF",X"FF",X"8F",X"F8",X"FF",X"FF",X"8F",X"F8",X"8F",X"FF",
		X"8F",X"F8",X"8F",X"FF",X"CF",X"F8",X"8F",X"FF",X"9F",X"F8",X"8F",X"FF",X"8F",X"F8",X"8F",X"FF",
		X"55",X"F9",X"99",X"99",X"55",X"FF",X"FF",X"FF",X"5F",X"F5",X"55",X"55",X"5F",X"75",X"55",X"55",
		X"55",X"F5",X"55",X"55",X"5F",X"75",X"55",X"55",X"55",X"F5",X"55",X"55",X"55",X"F5",X"55",X"55",
		X"FF",X"2F",X"FF",X"FF",X"F5",X"22",X"55",X"55",X"FF",X"7F",X"55",X"55",X"5F",X"F5",X"5F",X"5F",
		X"5F",X"F5",X"55",X"5F",X"FF",X"2F",X"55",X"5F",X"FF",X"72",X"5F",X"55",X"5F",X"F5",X"5F",X"55",
		X"A8",X"F5",X"8F",X"FF",X"88",X"F5",X"8F",X"FF",X"88",X"55",X"5F",X"FF",X"88",X"F5",X"8F",X"FF",
		X"88",X"F5",X"9F",X"FF",X"88",X"F8",X"9F",X"FF",X"88",X"58",X"95",X"F5",X"88",X"F5",X"85",X"5F",
		X"88",X"F5",X"85",X"F5",X"89",X"F9",X"8F",X"FF",X"99",X"F9",X"8F",X"FF",X"99",X"F9",X"8F",X"FF",
		X"99",X"DD",X"8F",X"FF",X"99",X"DD",X"8F",X"FF",X"99",X"DD",X"AF",X"FF",X"99",X"DD",X"AF",X"FF",
		X"CC",X"DD",X"AF",X"FF",X"AA",X"DD",X"AF",X"FF",X"EE",X"DD",X"AF",X"FF",X"79",X"DD",X"AF",X"FF",
		X"79",X"DD",X"AF",X"FF",X"79",X"DD",X"AF",X"FF",X"79",X"DD",X"AF",X"FF",X"79",X"DD",X"AF",X"FF",
		X"79",X"DD",X"AF",X"FF",X"79",X"DD",X"AF",X"FF",X"79",X"DD",X"AF",X"FF",X"79",X"DD",X"AF",X"FF",
		X"79",X"DD",X"AF",X"FF",X"79",X"DD",X"AF",X"FF",X"79",X"DD",X"AF",X"FF",X"79",X"DD",X"AF",X"FF",
		X"99",X"99",X"99",X"99",X"FF",X"FF",X"FF",X"77",X"55",X"55",X"55",X"77",X"55",X"5F",X"55",X"77",
		X"55",X"55",X"55",X"77",X"55",X"5F",X"55",X"F7",X"55",X"5F",X"55",X"5F",X"55",X"52",X"55",X"5F",
		X"FF",X"2F",X"FF",X"FF",X"F5",X"F5",X"5F",X"5F",X"55",X"F5",X"55",X"F7",X"55",X"F5",X"55",X"F7",
		X"55",X"F5",X"5F",X"5F",X"55",X"F5",X"55",X"F7",X"55",X"F5",X"5F",X"F7",X"55",X"F5",X"55",X"57",
		X"CF",X"22",X"22",X"77",X"7F",X"22",X"22",X"77",X"7F",X"22",X"CC",X"77",X"EF",X"22",X"CC",X"EE",
		X"AA",X"FF",X"FA",X"EE",X"FD",X"FF",X"F7",X"77",X"CD",X"AA",X"F7",X"C7",X"7D",X"EE",X"F7",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"FF",X"FF",X"FF",X"77",X"77",X"AA",X"A7",X"77",
		X"78",X"CC",X"A7",X"7F",X"78",X"CC",X"A7",X"7C",X"78",X"CC",X"A8",X"88",X"88",X"22",X"A8",X"88");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
